
//------> ./myproject_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module converterBlock_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./myproject_ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module converterBlock_ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./myproject.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
// 
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Sun Jan 15 03:49:02 2023
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core
// ------------------------------------------------------------------


module converterBlock_myproject_core (
  clk, rst, input_1_rsc_dat, layer7_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [95:0] input_1_rsc_dat;
  output [1:0] layer7_out_rsc_dat;
  input [4095:0] w2_rsc_dat;
  input [255:0] b2_rsc_dat;
  input [767:0] w5_rsc_dat;
  input [11:0] b5_rsc_dat;


  // Interconnect Declarations
  wire [95:0] input_1_rsci_idat;
  reg [1:0] layer7_out_rsci_idat;
  wire [4095:0] w2_rsci_idat;
  wire [255:0] b2_rsci_idat;
  wire [767:0] w5_rsci_idat;
  wire [11:0] b5_rsci_idat;
  wire [9:0] Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1;
  wire [15:0] nl_Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1;
  wire [7:0] Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1;
  wire [11:0] nl_Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1;
  wire [9:0] Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1;
  wire [15:0] nl_Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1;
  wire [9:0] Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1;
  wire [15:0] nl_Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire layer4_out_0_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_6_5;
  wire layer4_out_conc_4_7;
  wire [1:0] layer4_out_conc_4_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_6_5;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_7;
  wire [1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_6_5;
  wire [4:0] Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1;
  wire [4:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1;
  wire [4:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_8_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_8_1;

  wire[1:0] argmax_else_mux_nl;
  wire argmax_else_if_argmax_else_if_argmax_else_if_nor_nl;
  wire[10:0] argmax_else_aelse_acc_nl;
  wire[11:0] nl_argmax_else_aelse_acc_nl;
  wire[10:0] argmax_else_if_acc_nl;
  wire[11:0] nl_argmax_else_if_acc_nl;
  wire argmax_if_argmax_if_argmax_if_nor_nl;
  wire[10:0] argmax_aelse_acc_nl;
  wire[11:0] nl_argmax_aelse_acc_nl;
  wire[10:0] argmax_if_acc_nl;
  wire[11:0] nl_argmax_if_acc_nl;
  wire[7:0] Accum2_acc_946_nl;
  wire[8:0] nl_Accum2_acc_946_nl;
  wire[7:0] Product1_16_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_9_nl;
  wire[8:0] nl_Accum2_acc_9_nl;
  wire[7:0] Product1_16_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_16_nl;
  wire[8:0] nl_Accum2_acc_16_nl;
  wire[7:0] Product1_16_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_31_nl;
  wire[8:0] nl_Accum2_acc_31_nl;
  wire[7:0] Product1_16_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_46_nl;
  wire[8:0] nl_Accum2_acc_46_nl;
  wire[7:0] Product1_16_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_61_nl;
  wire[8:0] nl_Accum2_acc_61_nl;
  wire[7:0] Product1_16_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_76_nl;
  wire[8:0] nl_Accum2_acc_76_nl;
  wire[7:0] Product1_16_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_91_nl;
  wire[8:0] nl_Accum2_acc_91_nl;
  wire[7:0] Product1_16_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_106_nl;
  wire[8:0] nl_Accum2_acc_106_nl;
  wire[7:0] Product1_16_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_121_nl;
  wire[8:0] nl_Accum2_acc_121_nl;
  wire[7:0] Product1_16_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_136_nl;
  wire[8:0] nl_Accum2_acc_136_nl;
  wire[7:0] Product1_16_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_151_nl;
  wire[8:0] nl_Accum2_acc_151_nl;
  wire[7:0] Product1_16_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_166_nl;
  wire[8:0] nl_Accum2_acc_166_nl;
  wire[7:0] Product1_16_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_181_nl;
  wire[8:0] nl_Accum2_acc_181_nl;
  wire[7:0] Product1_16_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_196_nl;
  wire[8:0] nl_Accum2_acc_196_nl;
  wire[7:0] Product1_16_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_211_nl;
  wire[8:0] nl_Accum2_acc_211_nl;
  wire[7:0] Product1_16_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_226_nl;
  wire[8:0] nl_Accum2_acc_226_nl;
  wire[7:0] Product1_16_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_241_nl;
  wire[8:0] nl_Accum2_acc_241_nl;
  wire[7:0] Product1_16_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_256_nl;
  wire[8:0] nl_Accum2_acc_256_nl;
  wire[7:0] Product1_16_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_271_nl;
  wire[8:0] nl_Accum2_acc_271_nl;
  wire[7:0] Product1_16_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_286_nl;
  wire[8:0] nl_Accum2_acc_286_nl;
  wire[7:0] Product1_16_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_301_nl;
  wire[8:0] nl_Accum2_acc_301_nl;
  wire[7:0] Product1_16_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_316_nl;
  wire[8:0] nl_Accum2_acc_316_nl;
  wire[7:0] Product1_16_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_331_nl;
  wire[8:0] nl_Accum2_acc_331_nl;
  wire[7:0] Product1_16_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_346_nl;
  wire[8:0] nl_Accum2_acc_346_nl;
  wire[7:0] Product1_16_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_361_nl;
  wire[8:0] nl_Accum2_acc_361_nl;
  wire[7:0] Product1_16_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_376_nl;
  wire[8:0] nl_Accum2_acc_376_nl;
  wire[7:0] Product1_16_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_391_nl;
  wire[8:0] nl_Accum2_acc_391_nl;
  wire[7:0] Product1_16_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_406_nl;
  wire[8:0] nl_Accum2_acc_406_nl;
  wire[7:0] Product1_16_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_421_nl;
  wire[8:0] nl_Accum2_acc_421_nl;
  wire[7:0] Product1_16_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_436_nl;
  wire[8:0] nl_Accum2_acc_436_nl;
  wire[7:0] Product1_16_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_451_nl;
  wire[8:0] nl_Accum2_acc_451_nl;
  wire[7:0] Product1_16_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_466_nl;
  wire[8:0] nl_Accum2_acc_466_nl;
  wire[7:0] Product1_16_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_481_nl;
  wire[8:0] nl_Accum2_acc_481_nl;
  wire[7:0] Product1_16_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_496_nl;
  wire[8:0] nl_Accum2_acc_496_nl;
  wire[7:0] Product1_16_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_511_nl;
  wire[8:0] nl_Accum2_acc_511_nl;
  wire[7:0] Product1_16_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_526_nl;
  wire[8:0] nl_Accum2_acc_526_nl;
  wire[7:0] Product1_16_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_541_nl;
  wire[8:0] nl_Accum2_acc_541_nl;
  wire[7:0] Product1_16_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_556_nl;
  wire[8:0] nl_Accum2_acc_556_nl;
  wire[7:0] Product1_16_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_571_nl;
  wire[8:0] nl_Accum2_acc_571_nl;
  wire[7:0] Product1_16_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_586_nl;
  wire[8:0] nl_Accum2_acc_586_nl;
  wire[7:0] Product1_16_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_601_nl;
  wire[8:0] nl_Accum2_acc_601_nl;
  wire[7:0] Product1_16_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_616_nl;
  wire[8:0] nl_Accum2_acc_616_nl;
  wire[7:0] Product1_16_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_631_nl;
  wire[8:0] nl_Accum2_acc_631_nl;
  wire[7:0] Product1_16_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_646_nl;
  wire[8:0] nl_Accum2_acc_646_nl;
  wire[7:0] Product1_16_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_661_nl;
  wire[8:0] nl_Accum2_acc_661_nl;
  wire[7:0] Product1_16_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_676_nl;
  wire[8:0] nl_Accum2_acc_676_nl;
  wire[7:0] Product1_16_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_691_nl;
  wire[8:0] nl_Accum2_acc_691_nl;
  wire[7:0] Product1_16_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_706_nl;
  wire[8:0] nl_Accum2_acc_706_nl;
  wire[7:0] Product1_16_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_721_nl;
  wire[8:0] nl_Accum2_acc_721_nl;
  wire[7:0] Product1_16_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_736_nl;
  wire[8:0] nl_Accum2_acc_736_nl;
  wire[7:0] Product1_16_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_751_nl;
  wire[8:0] nl_Accum2_acc_751_nl;
  wire[7:0] Product1_16_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_766_nl;
  wire[8:0] nl_Accum2_acc_766_nl;
  wire[7:0] Product1_16_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_781_nl;
  wire[8:0] nl_Accum2_acc_781_nl;
  wire[7:0] Product1_16_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_796_nl;
  wire[8:0] nl_Accum2_acc_796_nl;
  wire[7:0] Product1_16_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_811_nl;
  wire[8:0] nl_Accum2_acc_811_nl;
  wire[7:0] Product1_16_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_826_nl;
  wire[8:0] nl_Accum2_acc_826_nl;
  wire[7:0] Product1_16_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_841_nl;
  wire[8:0] nl_Accum2_acc_841_nl;
  wire[7:0] Product1_16_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_856_nl;
  wire[8:0] nl_Accum2_acc_856_nl;
  wire[7:0] Product1_16_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_871_nl;
  wire[8:0] nl_Accum2_acc_871_nl;
  wire[7:0] Product1_16_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_886_nl;
  wire[8:0] nl_Accum2_acc_886_nl;
  wire[7:0] Product1_16_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_901_nl;
  wire[8:0] nl_Accum2_acc_901_nl;
  wire[7:0] Product1_16_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_916_nl;
  wire[8:0] nl_Accum2_acc_916_nl;
  wire[7:0] Product1_16_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Accum2_acc_931_nl;
  wire[8:0] nl_Accum2_acc_931_nl;
  wire[7:0] Product1_16_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_16_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_1_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_1_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_2_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_2_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_3_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_3_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_4_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_4_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_5_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_5_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_6_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_6_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_7_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_7_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_12_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_12_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_13_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_13_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_14_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_14_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_15_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_15_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_8_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_8_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_9_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_9_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_10_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_10_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[7:0] Product1_11_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [10:0] nl_Product1_11_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[9:0] Accum2_1_acc_127_nl;
  wire[14:0] nl_Accum2_1_acc_127_nl;
  wire[11:0] Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[4:0] Accum2_1_acc_192_nl;
  wire[5:0] nl_Accum2_1_acc_192_nl;
  wire[11:0] Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[9:0] Accum2_1_acc_190_nl;
  wire[14:0] nl_Accum2_1_acc_190_nl;
  wire[11:0] Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[4:0] Accum2_1_acc_193_nl;
  wire[5:0] nl_Accum2_1_acc_193_nl;
  wire[11:0] Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[9:0] Accum2_1_acc_nl;
  wire[14:0] nl_Accum2_1_acc_nl;
  wire[11:0] Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[4:0] Accum2_1_acc_191_nl;
  wire[5:0] nl_Accum2_1_acc_191_nl;
  wire[11:0] Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[11:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [12:0] nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[8:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl;
  wire[9:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;
  wire[1:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl;

  // Interconnect Declarations for Component Instantiations 
  converterBlock_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd96)) input_1_rsci (
      .dat(input_1_rsc_dat),
      .idat(input_1_rsci_idat)
    );
  converterBlock_ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd2)) layer7_out_rsci (
      .idat(layer7_out_rsci_idat),
      .dat(layer7_out_rsc_dat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd4096)) w2_rsci (
      .dat(w2_rsc_dat),
      .idat(w2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd256)) b2_rsci (
      .dat(b2_rsc_dat),
      .idat(b2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd768)) w5_rsci (
      .dat(w5_rsc_dat),
      .idat(w5_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd12)) b5_rsci (
      .dat(b5_rsc_dat),
      .idat(b5_rsci_idat)
    );
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1 = (Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3843:3840]));
  assign Product1_16_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_946_nl = Product1_16_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[3:0]);
  assign Accum2_acc_946_nl = nl_Accum2_acc_946_nl[7:0];
  assign nl_Product1_1_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[3:0]));
  assign Product1_1_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[259:256]));
  assign Product1_2_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[515:512]));
  assign Product1_3_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[771:768]));
  assign Product1_4_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1027:1024]));
  assign Product1_5_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1283:1280]));
  assign Product1_6_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1539:1536]));
  assign Product1_7_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2819:2816]));
  assign Product1_12_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3075:3072]));
  assign Product1_13_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3331:3328]));
  assign Product1_14_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3587:3584]));
  assign Product1_15_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1795:1792]));
  assign Product1_8_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2051:2048]));
  assign Product1_9_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2307:2304]));
  assign Product1_10_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2563:2560]));
  assign Product1_11_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1 = Accum2_acc_946_nl + Product1_1_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_1_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1 = nl_Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 = (Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3847:3844]));
  assign Product1_16_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_9_nl = Product1_16_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[7:4]);
  assign Accum2_acc_9_nl = nl_Accum2_acc_9_nl[7:0];
  assign nl_Product1_1_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[7:4]));
  assign Product1_1_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[263:260]));
  assign Product1_2_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[519:516]));
  assign Product1_3_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[775:772]));
  assign Product1_4_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1031:1028]));
  assign Product1_5_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1287:1284]));
  assign Product1_6_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1543:1540]));
  assign Product1_7_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2823:2820]));
  assign Product1_12_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3079:3076]));
  assign Product1_13_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3335:3332]));
  assign Product1_14_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3591:3588]));
  assign Product1_15_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1799:1796]));
  assign Product1_8_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2055:2052]));
  assign Product1_9_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2311:2308]));
  assign Product1_10_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2567:2564]));
  assign Product1_11_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1 = Accum2_acc_9_nl + Product1_1_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_2_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 = (Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3851:3848]));
  assign Product1_16_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_16_nl = Product1_16_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[11:8]);
  assign Accum2_acc_16_nl = nl_Accum2_acc_16_nl[7:0];
  assign nl_Product1_1_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[11:8]));
  assign Product1_1_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[267:264]));
  assign Product1_2_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[523:520]));
  assign Product1_3_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[779:776]));
  assign Product1_4_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1035:1032]));
  assign Product1_5_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1291:1288]));
  assign Product1_6_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1547:1544]));
  assign Product1_7_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2827:2824]));
  assign Product1_12_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3083:3080]));
  assign Product1_13_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3339:3336]));
  assign Product1_14_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3595:3592]));
  assign Product1_15_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1803:1800]));
  assign Product1_8_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2059:2056]));
  assign Product1_9_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2315:2312]));
  assign Product1_10_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2571:2568]));
  assign Product1_11_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1 = Accum2_acc_16_nl + Product1_1_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_3_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 = (Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3855:3852]));
  assign Product1_16_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_31_nl = Product1_16_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[15:12]);
  assign Accum2_acc_31_nl = nl_Accum2_acc_31_nl[7:0];
  assign nl_Product1_1_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[15:12]));
  assign Product1_1_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[271:268]));
  assign Product1_2_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[527:524]));
  assign Product1_3_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[783:780]));
  assign Product1_4_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1039:1036]));
  assign Product1_5_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1295:1292]));
  assign Product1_6_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1551:1548]));
  assign Product1_7_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2831:2828]));
  assign Product1_12_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3087:3084]));
  assign Product1_13_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3343:3340]));
  assign Product1_14_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3599:3596]));
  assign Product1_15_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1807:1804]));
  assign Product1_8_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2063:2060]));
  assign Product1_9_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2319:2316]));
  assign Product1_10_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2575:2572]));
  assign Product1_11_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1 = Accum2_acc_31_nl + Product1_1_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_4_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 = (Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3859:3856]));
  assign Product1_16_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_46_nl = Product1_16_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[19:16]);
  assign Accum2_acc_46_nl = nl_Accum2_acc_46_nl[7:0];
  assign nl_Product1_1_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[19:16]));
  assign Product1_1_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[275:272]));
  assign Product1_2_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[531:528]));
  assign Product1_3_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[787:784]));
  assign Product1_4_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1043:1040]));
  assign Product1_5_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1299:1296]));
  assign Product1_6_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1555:1552]));
  assign Product1_7_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2835:2832]));
  assign Product1_12_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3091:3088]));
  assign Product1_13_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3347:3344]));
  assign Product1_14_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3603:3600]));
  assign Product1_15_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1811:1808]));
  assign Product1_8_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2067:2064]));
  assign Product1_9_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2323:2320]));
  assign Product1_10_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2579:2576]));
  assign Product1_11_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1 = Accum2_acc_46_nl + Product1_1_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_5_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 = (Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3863:3860]));
  assign Product1_16_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_61_nl = Product1_16_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[23:20]);
  assign Accum2_acc_61_nl = nl_Accum2_acc_61_nl[7:0];
  assign nl_Product1_1_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[23:20]));
  assign Product1_1_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[279:276]));
  assign Product1_2_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[535:532]));
  assign Product1_3_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[791:788]));
  assign Product1_4_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1047:1044]));
  assign Product1_5_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1303:1300]));
  assign Product1_6_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1559:1556]));
  assign Product1_7_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2839:2836]));
  assign Product1_12_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3095:3092]));
  assign Product1_13_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3351:3348]));
  assign Product1_14_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3607:3604]));
  assign Product1_15_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1815:1812]));
  assign Product1_8_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2071:2068]));
  assign Product1_9_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2327:2324]));
  assign Product1_10_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2583:2580]));
  assign Product1_11_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1 = Accum2_acc_61_nl + Product1_1_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_6_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 = (Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3867:3864]));
  assign Product1_16_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_76_nl = Product1_16_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[27:24]);
  assign Accum2_acc_76_nl = nl_Accum2_acc_76_nl[7:0];
  assign nl_Product1_1_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[27:24]));
  assign Product1_1_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[283:280]));
  assign Product1_2_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[539:536]));
  assign Product1_3_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[795:792]));
  assign Product1_4_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1051:1048]));
  assign Product1_5_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1307:1304]));
  assign Product1_6_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1563:1560]));
  assign Product1_7_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2843:2840]));
  assign Product1_12_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3099:3096]));
  assign Product1_13_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3355:3352]));
  assign Product1_14_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3611:3608]));
  assign Product1_15_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1819:1816]));
  assign Product1_8_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2075:2072]));
  assign Product1_9_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2331:2328]));
  assign Product1_10_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2587:2584]));
  assign Product1_11_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1 = Accum2_acc_76_nl + Product1_1_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_7_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 = (Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3871:3868]));
  assign Product1_16_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_91_nl = Product1_16_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[31:28]);
  assign Accum2_acc_91_nl = nl_Accum2_acc_91_nl[7:0];
  assign nl_Product1_1_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[31:28]));
  assign Product1_1_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[287:284]));
  assign Product1_2_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[543:540]));
  assign Product1_3_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[799:796]));
  assign Product1_4_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1055:1052]));
  assign Product1_5_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1311:1308]));
  assign Product1_6_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1567:1564]));
  assign Product1_7_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2847:2844]));
  assign Product1_12_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3103:3100]));
  assign Product1_13_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3359:3356]));
  assign Product1_14_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3615:3612]));
  assign Product1_15_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1823:1820]));
  assign Product1_8_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2079:2076]));
  assign Product1_9_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2335:2332]));
  assign Product1_10_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2591:2588]));
  assign Product1_11_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1 = Accum2_acc_91_nl + Product1_1_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_8_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 = (Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3875:3872]));
  assign Product1_16_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_106_nl = Product1_16_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[35:32]);
  assign Accum2_acc_106_nl = nl_Accum2_acc_106_nl[7:0];
  assign nl_Product1_1_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[35:32]));
  assign Product1_1_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[291:288]));
  assign Product1_2_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[547:544]));
  assign Product1_3_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[803:800]));
  assign Product1_4_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1059:1056]));
  assign Product1_5_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1315:1312]));
  assign Product1_6_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1571:1568]));
  assign Product1_7_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2851:2848]));
  assign Product1_12_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3107:3104]));
  assign Product1_13_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3363:3360]));
  assign Product1_14_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3619:3616]));
  assign Product1_15_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1827:1824]));
  assign Product1_8_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2083:2080]));
  assign Product1_9_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2339:2336]));
  assign Product1_10_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2595:2592]));
  assign Product1_11_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1 = Accum2_acc_106_nl + Product1_1_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_3_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_4_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_5_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_6_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_9_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 = (Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3879:3876]));
  assign Product1_16_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_121_nl = Product1_16_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[39:36]);
  assign Accum2_acc_121_nl = nl_Accum2_acc_121_nl[7:0];
  assign nl_Product1_1_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[39:36]));
  assign Product1_1_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[295:292]));
  assign Product1_2_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[551:548]));
  assign Product1_3_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[807:804]));
  assign Product1_4_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1063:1060]));
  assign Product1_5_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1319:1316]));
  assign Product1_6_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1575:1572]));
  assign Product1_7_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2855:2852]));
  assign Product1_12_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3111:3108]));
  assign Product1_13_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3367:3364]));
  assign Product1_14_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3623:3620]));
  assign Product1_15_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1831:1828]));
  assign Product1_8_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2087:2084]));
  assign Product1_9_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2343:2340]));
  assign Product1_10_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2599:2596]));
  assign Product1_11_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1 = Accum2_acc_121_nl + Product1_1_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_10_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 = (Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3883:3880]));
  assign Product1_16_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_136_nl = Product1_16_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[43:40]);
  assign Accum2_acc_136_nl = nl_Accum2_acc_136_nl[7:0];
  assign nl_Product1_1_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[43:40]));
  assign Product1_1_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[299:296]));
  assign Product1_2_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[555:552]));
  assign Product1_3_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[811:808]));
  assign Product1_4_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1067:1064]));
  assign Product1_5_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1323:1320]));
  assign Product1_6_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1579:1576]));
  assign Product1_7_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2859:2856]));
  assign Product1_12_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3115:3112]));
  assign Product1_13_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3371:3368]));
  assign Product1_14_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3627:3624]));
  assign Product1_15_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1835:1832]));
  assign Product1_8_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2091:2088]));
  assign Product1_9_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2347:2344]));
  assign Product1_10_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2603:2600]));
  assign Product1_11_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1 = Accum2_acc_136_nl + Product1_1_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_11_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 = (Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3887:3884]));
  assign Product1_16_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_151_nl = Product1_16_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[47:44]);
  assign Accum2_acc_151_nl = nl_Accum2_acc_151_nl[7:0];
  assign nl_Product1_1_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[47:44]));
  assign Product1_1_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[303:300]));
  assign Product1_2_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[559:556]));
  assign Product1_3_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[815:812]));
  assign Product1_4_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1071:1068]));
  assign Product1_5_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1327:1324]));
  assign Product1_6_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1583:1580]));
  assign Product1_7_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2863:2860]));
  assign Product1_12_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3119:3116]));
  assign Product1_13_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3375:3372]));
  assign Product1_14_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3631:3628]));
  assign Product1_15_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1839:1836]));
  assign Product1_8_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2095:2092]));
  assign Product1_9_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2351:2348]));
  assign Product1_10_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2607:2604]));
  assign Product1_11_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1 = Accum2_acc_151_nl + Product1_1_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_12_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 = (Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3891:3888]));
  assign Product1_16_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_166_nl = Product1_16_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[51:48]);
  assign Accum2_acc_166_nl = nl_Accum2_acc_166_nl[7:0];
  assign nl_Product1_1_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[51:48]));
  assign Product1_1_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[307:304]));
  assign Product1_2_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[563:560]));
  assign Product1_3_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[819:816]));
  assign Product1_4_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1075:1072]));
  assign Product1_5_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1331:1328]));
  assign Product1_6_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1587:1584]));
  assign Product1_7_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2867:2864]));
  assign Product1_12_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3123:3120]));
  assign Product1_13_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3379:3376]));
  assign Product1_14_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3635:3632]));
  assign Product1_15_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1843:1840]));
  assign Product1_8_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2099:2096]));
  assign Product1_9_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2355:2352]));
  assign Product1_10_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2611:2608]));
  assign Product1_11_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1 = Accum2_acc_166_nl + Product1_1_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_13_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 = (Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3895:3892]));
  assign Product1_16_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_181_nl = Product1_16_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[55:52]);
  assign Accum2_acc_181_nl = nl_Accum2_acc_181_nl[7:0];
  assign nl_Product1_1_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[55:52]));
  assign Product1_1_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[311:308]));
  assign Product1_2_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[567:564]));
  assign Product1_3_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[823:820]));
  assign Product1_4_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1079:1076]));
  assign Product1_5_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1335:1332]));
  assign Product1_6_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1591:1588]));
  assign Product1_7_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2871:2868]));
  assign Product1_12_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3127:3124]));
  assign Product1_13_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3383:3380]));
  assign Product1_14_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3639:3636]));
  assign Product1_15_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1847:1844]));
  assign Product1_8_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2103:2100]));
  assign Product1_9_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2359:2356]));
  assign Product1_10_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2615:2612]));
  assign Product1_11_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1 = Accum2_acc_181_nl + Product1_1_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_14_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 = (Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3899:3896]));
  assign Product1_16_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_196_nl = Product1_16_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[59:56]);
  assign Accum2_acc_196_nl = nl_Accum2_acc_196_nl[7:0];
  assign nl_Product1_1_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[59:56]));
  assign Product1_1_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[315:312]));
  assign Product1_2_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[571:568]));
  assign Product1_3_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[827:824]));
  assign Product1_4_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1083:1080]));
  assign Product1_5_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1339:1336]));
  assign Product1_6_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1595:1592]));
  assign Product1_7_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2875:2872]));
  assign Product1_12_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3131:3128]));
  assign Product1_13_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3387:3384]));
  assign Product1_14_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3643:3640]));
  assign Product1_15_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1851:1848]));
  assign Product1_8_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2107:2104]));
  assign Product1_9_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2363:2360]));
  assign Product1_10_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2619:2616]));
  assign Product1_11_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1 = Accum2_acc_196_nl + Product1_1_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_15_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 = (Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3903:3900]));
  assign Product1_16_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_211_nl = Product1_16_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[63:60]);
  assign Accum2_acc_211_nl = nl_Accum2_acc_211_nl[7:0];
  assign nl_Product1_1_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[63:60]));
  assign Product1_1_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[319:316]));
  assign Product1_2_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[575:572]));
  assign Product1_3_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[831:828]));
  assign Product1_4_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1087:1084]));
  assign Product1_5_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1343:1340]));
  assign Product1_6_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1599:1596]));
  assign Product1_7_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2879:2876]));
  assign Product1_12_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3135:3132]));
  assign Product1_13_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3391:3388]));
  assign Product1_14_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3647:3644]));
  assign Product1_15_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1855:1852]));
  assign Product1_8_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2111:2108]));
  assign Product1_9_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2367:2364]));
  assign Product1_10_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2623:2620]));
  assign Product1_11_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1 = Accum2_acc_211_nl + Product1_1_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_16_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 = (Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3907:3904]));
  assign Product1_16_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_226_nl = Product1_16_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[67:64]);
  assign Accum2_acc_226_nl = nl_Accum2_acc_226_nl[7:0];
  assign nl_Product1_1_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[67:64]));
  assign Product1_1_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[323:320]));
  assign Product1_2_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[579:576]));
  assign Product1_3_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[835:832]));
  assign Product1_4_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1091:1088]));
  assign Product1_5_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1347:1344]));
  assign Product1_6_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1603:1600]));
  assign Product1_7_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2883:2880]));
  assign Product1_12_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3139:3136]));
  assign Product1_13_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3395:3392]));
  assign Product1_14_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3651:3648]));
  assign Product1_15_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1859:1856]));
  assign Product1_8_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2115:2112]));
  assign Product1_9_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2371:2368]));
  assign Product1_10_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2627:2624]));
  assign Product1_11_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1 = Accum2_acc_226_nl + Product1_1_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_17_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 = (Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3911:3908]));
  assign Product1_16_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_241_nl = Product1_16_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[71:68]);
  assign Accum2_acc_241_nl = nl_Accum2_acc_241_nl[7:0];
  assign nl_Product1_1_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[71:68]));
  assign Product1_1_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[327:324]));
  assign Product1_2_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[583:580]));
  assign Product1_3_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[839:836]));
  assign Product1_4_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1095:1092]));
  assign Product1_5_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1351:1348]));
  assign Product1_6_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1607:1604]));
  assign Product1_7_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2887:2884]));
  assign Product1_12_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3143:3140]));
  assign Product1_13_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3399:3396]));
  assign Product1_14_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3655:3652]));
  assign Product1_15_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1863:1860]));
  assign Product1_8_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2119:2116]));
  assign Product1_9_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2375:2372]));
  assign Product1_10_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2631:2628]));
  assign Product1_11_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1 = Accum2_acc_241_nl + Product1_1_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_18_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 = (Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3915:3912]));
  assign Product1_16_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_256_nl = Product1_16_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[75:72]);
  assign Accum2_acc_256_nl = nl_Accum2_acc_256_nl[7:0];
  assign nl_Product1_1_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[75:72]));
  assign Product1_1_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[331:328]));
  assign Product1_2_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[587:584]));
  assign Product1_3_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[843:840]));
  assign Product1_4_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1099:1096]));
  assign Product1_5_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1355:1352]));
  assign Product1_6_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1611:1608]));
  assign Product1_7_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2891:2888]));
  assign Product1_12_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3147:3144]));
  assign Product1_13_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3403:3400]));
  assign Product1_14_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3659:3656]));
  assign Product1_15_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1867:1864]));
  assign Product1_8_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2123:2120]));
  assign Product1_9_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2379:2376]));
  assign Product1_10_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2635:2632]));
  assign Product1_11_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1 = Accum2_acc_256_nl + Product1_1_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_19_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 = (Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3919:3916]));
  assign Product1_16_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_271_nl = Product1_16_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[79:76]);
  assign Accum2_acc_271_nl = nl_Accum2_acc_271_nl[7:0];
  assign nl_Product1_1_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[79:76]));
  assign Product1_1_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[335:332]));
  assign Product1_2_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[591:588]));
  assign Product1_3_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[847:844]));
  assign Product1_4_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1103:1100]));
  assign Product1_5_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1359:1356]));
  assign Product1_6_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1615:1612]));
  assign Product1_7_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2895:2892]));
  assign Product1_12_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3151:3148]));
  assign Product1_13_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3407:3404]));
  assign Product1_14_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3663:3660]));
  assign Product1_15_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1871:1868]));
  assign Product1_8_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2127:2124]));
  assign Product1_9_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2383:2380]));
  assign Product1_10_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2639:2636]));
  assign Product1_11_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1 = Accum2_acc_271_nl + Product1_1_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_20_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 = (Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3923:3920]));
  assign Product1_16_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_286_nl = Product1_16_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[83:80]);
  assign Accum2_acc_286_nl = nl_Accum2_acc_286_nl[7:0];
  assign nl_Product1_1_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[83:80]));
  assign Product1_1_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[339:336]));
  assign Product1_2_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[595:592]));
  assign Product1_3_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[851:848]));
  assign Product1_4_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1107:1104]));
  assign Product1_5_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1363:1360]));
  assign Product1_6_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1619:1616]));
  assign Product1_7_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2899:2896]));
  assign Product1_12_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3155:3152]));
  assign Product1_13_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3411:3408]));
  assign Product1_14_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3667:3664]));
  assign Product1_15_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1875:1872]));
  assign Product1_8_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2131:2128]));
  assign Product1_9_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2387:2384]));
  assign Product1_10_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2643:2640]));
  assign Product1_11_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1 = Accum2_acc_286_nl + Product1_1_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_21_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 = (Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3927:3924]));
  assign Product1_16_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_301_nl = Product1_16_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[87:84]);
  assign Accum2_acc_301_nl = nl_Accum2_acc_301_nl[7:0];
  assign nl_Product1_1_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[87:84]));
  assign Product1_1_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[343:340]));
  assign Product1_2_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[599:596]));
  assign Product1_3_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[855:852]));
  assign Product1_4_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1111:1108]));
  assign Product1_5_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1367:1364]));
  assign Product1_6_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1623:1620]));
  assign Product1_7_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2903:2900]));
  assign Product1_12_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3159:3156]));
  assign Product1_13_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3415:3412]));
  assign Product1_14_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3671:3668]));
  assign Product1_15_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1879:1876]));
  assign Product1_8_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2135:2132]));
  assign Product1_9_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2391:2388]));
  assign Product1_10_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2647:2644]));
  assign Product1_11_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1 = Accum2_acc_301_nl + Product1_1_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_22_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 = (Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3931:3928]));
  assign Product1_16_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_316_nl = Product1_16_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[91:88]);
  assign Accum2_acc_316_nl = nl_Accum2_acc_316_nl[7:0];
  assign nl_Product1_1_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[91:88]));
  assign Product1_1_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[347:344]));
  assign Product1_2_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[603:600]));
  assign Product1_3_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[859:856]));
  assign Product1_4_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1115:1112]));
  assign Product1_5_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1371:1368]));
  assign Product1_6_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1627:1624]));
  assign Product1_7_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2907:2904]));
  assign Product1_12_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3163:3160]));
  assign Product1_13_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3419:3416]));
  assign Product1_14_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3675:3672]));
  assign Product1_15_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1883:1880]));
  assign Product1_8_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2139:2136]));
  assign Product1_9_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2395:2392]));
  assign Product1_10_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2651:2648]));
  assign Product1_11_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1 = Accum2_acc_316_nl + Product1_1_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_23_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 = (Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3935:3932]));
  assign Product1_16_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_331_nl = Product1_16_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[95:92]);
  assign Accum2_acc_331_nl = nl_Accum2_acc_331_nl[7:0];
  assign nl_Product1_1_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[95:92]));
  assign Product1_1_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[351:348]));
  assign Product1_2_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[607:604]));
  assign Product1_3_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[863:860]));
  assign Product1_4_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1119:1116]));
  assign Product1_5_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1375:1372]));
  assign Product1_6_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1631:1628]));
  assign Product1_7_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2911:2908]));
  assign Product1_12_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3167:3164]));
  assign Product1_13_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3423:3420]));
  assign Product1_14_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3679:3676]));
  assign Product1_15_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1887:1884]));
  assign Product1_8_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2143:2140]));
  assign Product1_9_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2399:2396]));
  assign Product1_10_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2655:2652]));
  assign Product1_11_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1 = Accum2_acc_331_nl + Product1_1_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_24_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 = (Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3939:3936]));
  assign Product1_16_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_346_nl = Product1_16_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[99:96]);
  assign Accum2_acc_346_nl = nl_Accum2_acc_346_nl[7:0];
  assign nl_Product1_1_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[99:96]));
  assign Product1_1_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[355:352]));
  assign Product1_2_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[611:608]));
  assign Product1_3_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[867:864]));
  assign Product1_4_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1123:1120]));
  assign Product1_5_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1379:1376]));
  assign Product1_6_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1635:1632]));
  assign Product1_7_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2915:2912]));
  assign Product1_12_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3171:3168]));
  assign Product1_13_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3427:3424]));
  assign Product1_14_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3683:3680]));
  assign Product1_15_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1891:1888]));
  assign Product1_8_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2147:2144]));
  assign Product1_9_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2403:2400]));
  assign Product1_10_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2659:2656]));
  assign Product1_11_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1 = Accum2_acc_346_nl + Product1_1_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_25_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 = (Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3943:3940]));
  assign Product1_16_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_361_nl = Product1_16_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[103:100]);
  assign Accum2_acc_361_nl = nl_Accum2_acc_361_nl[7:0];
  assign nl_Product1_1_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[103:100]));
  assign Product1_1_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[359:356]));
  assign Product1_2_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[615:612]));
  assign Product1_3_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[871:868]));
  assign Product1_4_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1127:1124]));
  assign Product1_5_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1383:1380]));
  assign Product1_6_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1639:1636]));
  assign Product1_7_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2919:2916]));
  assign Product1_12_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3175:3172]));
  assign Product1_13_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3431:3428]));
  assign Product1_14_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3687:3684]));
  assign Product1_15_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1895:1892]));
  assign Product1_8_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2151:2148]));
  assign Product1_9_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2407:2404]));
  assign Product1_10_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2663:2660]));
  assign Product1_11_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1 = Accum2_acc_361_nl + Product1_1_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_26_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 = (Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3947:3944]));
  assign Product1_16_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_376_nl = Product1_16_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[107:104]);
  assign Accum2_acc_376_nl = nl_Accum2_acc_376_nl[7:0];
  assign nl_Product1_1_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[107:104]));
  assign Product1_1_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[363:360]));
  assign Product1_2_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[619:616]));
  assign Product1_3_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[875:872]));
  assign Product1_4_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1131:1128]));
  assign Product1_5_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1387:1384]));
  assign Product1_6_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1643:1640]));
  assign Product1_7_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2923:2920]));
  assign Product1_12_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3179:3176]));
  assign Product1_13_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3435:3432]));
  assign Product1_14_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3691:3688]));
  assign Product1_15_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1899:1896]));
  assign Product1_8_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2155:2152]));
  assign Product1_9_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2411:2408]));
  assign Product1_10_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2667:2664]));
  assign Product1_11_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1 = Accum2_acc_376_nl + Product1_1_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_27_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 = (Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3951:3948]));
  assign Product1_16_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_391_nl = Product1_16_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[111:108]);
  assign Accum2_acc_391_nl = nl_Accum2_acc_391_nl[7:0];
  assign nl_Product1_1_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[111:108]));
  assign Product1_1_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[367:364]));
  assign Product1_2_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[623:620]));
  assign Product1_3_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[879:876]));
  assign Product1_4_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1135:1132]));
  assign Product1_5_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1391:1388]));
  assign Product1_6_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1647:1644]));
  assign Product1_7_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2927:2924]));
  assign Product1_12_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3183:3180]));
  assign Product1_13_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3439:3436]));
  assign Product1_14_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3695:3692]));
  assign Product1_15_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1903:1900]));
  assign Product1_8_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2159:2156]));
  assign Product1_9_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2415:2412]));
  assign Product1_10_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2671:2668]));
  assign Product1_11_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1 = Accum2_acc_391_nl + Product1_1_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_28_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 = (Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3955:3952]));
  assign Product1_16_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_406_nl = Product1_16_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[115:112]);
  assign Accum2_acc_406_nl = nl_Accum2_acc_406_nl[7:0];
  assign nl_Product1_1_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[115:112]));
  assign Product1_1_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[371:368]));
  assign Product1_2_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[627:624]));
  assign Product1_3_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[883:880]));
  assign Product1_4_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1139:1136]));
  assign Product1_5_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1395:1392]));
  assign Product1_6_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1651:1648]));
  assign Product1_7_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2931:2928]));
  assign Product1_12_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3187:3184]));
  assign Product1_13_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3443:3440]));
  assign Product1_14_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3699:3696]));
  assign Product1_15_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1907:1904]));
  assign Product1_8_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2163:2160]));
  assign Product1_9_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2419:2416]));
  assign Product1_10_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2675:2672]));
  assign Product1_11_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1 = Accum2_acc_406_nl + Product1_1_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_29_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 = (Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3959:3956]));
  assign Product1_16_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_421_nl = Product1_16_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[119:116]);
  assign Accum2_acc_421_nl = nl_Accum2_acc_421_nl[7:0];
  assign nl_Product1_1_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[119:116]));
  assign Product1_1_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[375:372]));
  assign Product1_2_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[631:628]));
  assign Product1_3_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[887:884]));
  assign Product1_4_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1143:1140]));
  assign Product1_5_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1399:1396]));
  assign Product1_6_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1655:1652]));
  assign Product1_7_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2935:2932]));
  assign Product1_12_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3191:3188]));
  assign Product1_13_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3447:3444]));
  assign Product1_14_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3703:3700]));
  assign Product1_15_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1911:1908]));
  assign Product1_8_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2167:2164]));
  assign Product1_9_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2423:2420]));
  assign Product1_10_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2679:2676]));
  assign Product1_11_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1 = Accum2_acc_421_nl + Product1_1_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_30_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 = (Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3963:3960]));
  assign Product1_16_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_436_nl = Product1_16_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[123:120]);
  assign Accum2_acc_436_nl = nl_Accum2_acc_436_nl[7:0];
  assign nl_Product1_1_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[123:120]));
  assign Product1_1_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[379:376]));
  assign Product1_2_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[635:632]));
  assign Product1_3_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[891:888]));
  assign Product1_4_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1147:1144]));
  assign Product1_5_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1403:1400]));
  assign Product1_6_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1659:1656]));
  assign Product1_7_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2939:2936]));
  assign Product1_12_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3195:3192]));
  assign Product1_13_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3451:3448]));
  assign Product1_14_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3707:3704]));
  assign Product1_15_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1915:1912]));
  assign Product1_8_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2171:2168]));
  assign Product1_9_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2427:2424]));
  assign Product1_10_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2683:2680]));
  assign Product1_11_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1 = Accum2_acc_436_nl + Product1_1_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_31_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 = (Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3967:3964]));
  assign Product1_16_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_451_nl = Product1_16_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[127:124]);
  assign Accum2_acc_451_nl = nl_Accum2_acc_451_nl[7:0];
  assign nl_Product1_1_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[127:124]));
  assign Product1_1_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[383:380]));
  assign Product1_2_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[639:636]));
  assign Product1_3_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[895:892]));
  assign Product1_4_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1151:1148]));
  assign Product1_5_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1407:1404]));
  assign Product1_6_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1663:1660]));
  assign Product1_7_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2943:2940]));
  assign Product1_12_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3199:3196]));
  assign Product1_13_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3455:3452]));
  assign Product1_14_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3711:3708]));
  assign Product1_15_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1919:1916]));
  assign Product1_8_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2175:2172]));
  assign Product1_9_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2431:2428]));
  assign Product1_10_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2687:2684]));
  assign Product1_11_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1 = Accum2_acc_451_nl + Product1_1_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_32_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 = (Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3971:3968]));
  assign Product1_16_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_466_nl = Product1_16_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[131:128]);
  assign Accum2_acc_466_nl = nl_Accum2_acc_466_nl[7:0];
  assign nl_Product1_1_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[131:128]));
  assign Product1_1_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[387:384]));
  assign Product1_2_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[643:640]));
  assign Product1_3_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[899:896]));
  assign Product1_4_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1155:1152]));
  assign Product1_5_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1411:1408]));
  assign Product1_6_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1667:1664]));
  assign Product1_7_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2947:2944]));
  assign Product1_12_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3203:3200]));
  assign Product1_13_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3459:3456]));
  assign Product1_14_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3715:3712]));
  assign Product1_15_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1923:1920]));
  assign Product1_8_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2179:2176]));
  assign Product1_9_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2435:2432]));
  assign Product1_10_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2691:2688]));
  assign Product1_11_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1 = Accum2_acc_466_nl + Product1_1_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_33_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 = (Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3975:3972]));
  assign Product1_16_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_481_nl = Product1_16_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[135:132]);
  assign Accum2_acc_481_nl = nl_Accum2_acc_481_nl[7:0];
  assign nl_Product1_1_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[135:132]));
  assign Product1_1_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[391:388]));
  assign Product1_2_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[647:644]));
  assign Product1_3_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[903:900]));
  assign Product1_4_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1159:1156]));
  assign Product1_5_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1415:1412]));
  assign Product1_6_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1671:1668]));
  assign Product1_7_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2951:2948]));
  assign Product1_12_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3207:3204]));
  assign Product1_13_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3463:3460]));
  assign Product1_14_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3719:3716]));
  assign Product1_15_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1927:1924]));
  assign Product1_8_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2183:2180]));
  assign Product1_9_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2439:2436]));
  assign Product1_10_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2695:2692]));
  assign Product1_11_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1 = Accum2_acc_481_nl + Product1_1_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_34_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 = (Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3979:3976]));
  assign Product1_16_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_496_nl = Product1_16_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[139:136]);
  assign Accum2_acc_496_nl = nl_Accum2_acc_496_nl[7:0];
  assign nl_Product1_1_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[139:136]));
  assign Product1_1_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[395:392]));
  assign Product1_2_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[651:648]));
  assign Product1_3_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[907:904]));
  assign Product1_4_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1163:1160]));
  assign Product1_5_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1419:1416]));
  assign Product1_6_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1675:1672]));
  assign Product1_7_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2955:2952]));
  assign Product1_12_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3211:3208]));
  assign Product1_13_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3467:3464]));
  assign Product1_14_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3723:3720]));
  assign Product1_15_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1931:1928]));
  assign Product1_8_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2187:2184]));
  assign Product1_9_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2443:2440]));
  assign Product1_10_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2699:2696]));
  assign Product1_11_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1 = Accum2_acc_496_nl + Product1_1_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_35_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 = (Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3983:3980]));
  assign Product1_16_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_511_nl = Product1_16_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[143:140]);
  assign Accum2_acc_511_nl = nl_Accum2_acc_511_nl[7:0];
  assign nl_Product1_1_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[143:140]));
  assign Product1_1_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[399:396]));
  assign Product1_2_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[655:652]));
  assign Product1_3_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[911:908]));
  assign Product1_4_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1167:1164]));
  assign Product1_5_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1423:1420]));
  assign Product1_6_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1679:1676]));
  assign Product1_7_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2959:2956]));
  assign Product1_12_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3215:3212]));
  assign Product1_13_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3471:3468]));
  assign Product1_14_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3727:3724]));
  assign Product1_15_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1935:1932]));
  assign Product1_8_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2191:2188]));
  assign Product1_9_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2447:2444]));
  assign Product1_10_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2703:2700]));
  assign Product1_11_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1 = Accum2_acc_511_nl + Product1_1_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_36_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 = (Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3987:3984]));
  assign Product1_16_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_526_nl = Product1_16_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[147:144]);
  assign Accum2_acc_526_nl = nl_Accum2_acc_526_nl[7:0];
  assign nl_Product1_1_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[147:144]));
  assign Product1_1_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[403:400]));
  assign Product1_2_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[659:656]));
  assign Product1_3_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[915:912]));
  assign Product1_4_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1171:1168]));
  assign Product1_5_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1427:1424]));
  assign Product1_6_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1683:1680]));
  assign Product1_7_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2963:2960]));
  assign Product1_12_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3219:3216]));
  assign Product1_13_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3475:3472]));
  assign Product1_14_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3731:3728]));
  assign Product1_15_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1939:1936]));
  assign Product1_8_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2195:2192]));
  assign Product1_9_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2451:2448]));
  assign Product1_10_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2707:2704]));
  assign Product1_11_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1 = Accum2_acc_526_nl + Product1_1_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_37_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 = (Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3991:3988]));
  assign Product1_16_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_541_nl = Product1_16_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[151:148]);
  assign Accum2_acc_541_nl = nl_Accum2_acc_541_nl[7:0];
  assign nl_Product1_1_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[151:148]));
  assign Product1_1_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[407:404]));
  assign Product1_2_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[663:660]));
  assign Product1_3_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[919:916]));
  assign Product1_4_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1175:1172]));
  assign Product1_5_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1431:1428]));
  assign Product1_6_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1687:1684]));
  assign Product1_7_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2967:2964]));
  assign Product1_12_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3223:3220]));
  assign Product1_13_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3479:3476]));
  assign Product1_14_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3735:3732]));
  assign Product1_15_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1943:1940]));
  assign Product1_8_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2199:2196]));
  assign Product1_9_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2455:2452]));
  assign Product1_10_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2711:2708]));
  assign Product1_11_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1 = Accum2_acc_541_nl + Product1_1_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_38_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 = (Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3995:3992]));
  assign Product1_16_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_556_nl = Product1_16_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[155:152]);
  assign Accum2_acc_556_nl = nl_Accum2_acc_556_nl[7:0];
  assign nl_Product1_1_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[155:152]));
  assign Product1_1_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[411:408]));
  assign Product1_2_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[667:664]));
  assign Product1_3_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[923:920]));
  assign Product1_4_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1179:1176]));
  assign Product1_5_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1435:1432]));
  assign Product1_6_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1691:1688]));
  assign Product1_7_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2971:2968]));
  assign Product1_12_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3227:3224]));
  assign Product1_13_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3483:3480]));
  assign Product1_14_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3739:3736]));
  assign Product1_15_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1947:1944]));
  assign Product1_8_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2203:2200]));
  assign Product1_9_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2459:2456]));
  assign Product1_10_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2715:2712]));
  assign Product1_11_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1 = Accum2_acc_556_nl + Product1_1_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_39_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 = (Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[3999:3996]));
  assign Product1_16_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_571_nl = Product1_16_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[159:156]);
  assign Accum2_acc_571_nl = nl_Accum2_acc_571_nl[7:0];
  assign nl_Product1_1_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[159:156]));
  assign Product1_1_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[415:412]));
  assign Product1_2_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[671:668]));
  assign Product1_3_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[927:924]));
  assign Product1_4_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1183:1180]));
  assign Product1_5_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1439:1436]));
  assign Product1_6_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1695:1692]));
  assign Product1_7_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2975:2972]));
  assign Product1_12_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3231:3228]));
  assign Product1_13_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3487:3484]));
  assign Product1_14_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3743:3740]));
  assign Product1_15_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1951:1948]));
  assign Product1_8_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2207:2204]));
  assign Product1_9_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2463:2460]));
  assign Product1_10_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2719:2716]));
  assign Product1_11_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1 = Accum2_acc_571_nl + Product1_1_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_40_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 = (Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4003:4000]));
  assign Product1_16_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_586_nl = Product1_16_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[163:160]);
  assign Accum2_acc_586_nl = nl_Accum2_acc_586_nl[7:0];
  assign nl_Product1_1_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[163:160]));
  assign Product1_1_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[419:416]));
  assign Product1_2_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[675:672]));
  assign Product1_3_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[931:928]));
  assign Product1_4_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1187:1184]));
  assign Product1_5_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1443:1440]));
  assign Product1_6_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1699:1696]));
  assign Product1_7_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2979:2976]));
  assign Product1_12_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3235:3232]));
  assign Product1_13_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3491:3488]));
  assign Product1_14_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3747:3744]));
  assign Product1_15_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1955:1952]));
  assign Product1_8_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2211:2208]));
  assign Product1_9_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2467:2464]));
  assign Product1_10_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2723:2720]));
  assign Product1_11_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1 = Accum2_acc_586_nl + Product1_1_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_41_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 = (Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4007:4004]));
  assign Product1_16_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_601_nl = Product1_16_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[167:164]);
  assign Accum2_acc_601_nl = nl_Accum2_acc_601_nl[7:0];
  assign nl_Product1_1_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[167:164]));
  assign Product1_1_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[423:420]));
  assign Product1_2_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[679:676]));
  assign Product1_3_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[935:932]));
  assign Product1_4_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1191:1188]));
  assign Product1_5_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1447:1444]));
  assign Product1_6_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1703:1700]));
  assign Product1_7_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2983:2980]));
  assign Product1_12_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3239:3236]));
  assign Product1_13_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3495:3492]));
  assign Product1_14_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3751:3748]));
  assign Product1_15_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1959:1956]));
  assign Product1_8_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2215:2212]));
  assign Product1_9_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2471:2468]));
  assign Product1_10_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2727:2724]));
  assign Product1_11_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1 = Accum2_acc_601_nl + Product1_1_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_42_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 = (Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4011:4008]));
  assign Product1_16_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_616_nl = Product1_16_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[171:168]);
  assign Accum2_acc_616_nl = nl_Accum2_acc_616_nl[7:0];
  assign nl_Product1_1_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[171:168]));
  assign Product1_1_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[427:424]));
  assign Product1_2_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[683:680]));
  assign Product1_3_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[939:936]));
  assign Product1_4_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1195:1192]));
  assign Product1_5_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1451:1448]));
  assign Product1_6_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1707:1704]));
  assign Product1_7_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2987:2984]));
  assign Product1_12_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3243:3240]));
  assign Product1_13_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3499:3496]));
  assign Product1_14_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3755:3752]));
  assign Product1_15_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1963:1960]));
  assign Product1_8_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2219:2216]));
  assign Product1_9_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2475:2472]));
  assign Product1_10_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2731:2728]));
  assign Product1_11_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1 = Accum2_acc_616_nl + Product1_1_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_43_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 = (Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4015:4012]));
  assign Product1_16_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_631_nl = Product1_16_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[175:172]);
  assign Accum2_acc_631_nl = nl_Accum2_acc_631_nl[7:0];
  assign nl_Product1_1_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[175:172]));
  assign Product1_1_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[431:428]));
  assign Product1_2_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[687:684]));
  assign Product1_3_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[943:940]));
  assign Product1_4_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1199:1196]));
  assign Product1_5_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1455:1452]));
  assign Product1_6_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1711:1708]));
  assign Product1_7_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2991:2988]));
  assign Product1_12_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3247:3244]));
  assign Product1_13_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3503:3500]));
  assign Product1_14_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3759:3756]));
  assign Product1_15_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1967:1964]));
  assign Product1_8_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2223:2220]));
  assign Product1_9_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2479:2476]));
  assign Product1_10_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2735:2732]));
  assign Product1_11_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1 = Accum2_acc_631_nl + Product1_1_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_44_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 = (Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4019:4016]));
  assign Product1_16_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_646_nl = Product1_16_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[179:176]);
  assign Accum2_acc_646_nl = nl_Accum2_acc_646_nl[7:0];
  assign nl_Product1_1_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[179:176]));
  assign Product1_1_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[435:432]));
  assign Product1_2_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[691:688]));
  assign Product1_3_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[947:944]));
  assign Product1_4_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1203:1200]));
  assign Product1_5_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1459:1456]));
  assign Product1_6_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1715:1712]));
  assign Product1_7_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2995:2992]));
  assign Product1_12_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3251:3248]));
  assign Product1_13_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3507:3504]));
  assign Product1_14_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3763:3760]));
  assign Product1_15_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1971:1968]));
  assign Product1_8_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2227:2224]));
  assign Product1_9_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2483:2480]));
  assign Product1_10_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2739:2736]));
  assign Product1_11_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1 = Accum2_acc_646_nl + Product1_1_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_45_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 = (Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4023:4020]));
  assign Product1_16_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_661_nl = Product1_16_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[183:180]);
  assign Accum2_acc_661_nl = nl_Accum2_acc_661_nl[7:0];
  assign nl_Product1_1_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[183:180]));
  assign Product1_1_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[439:436]));
  assign Product1_2_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[695:692]));
  assign Product1_3_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[951:948]));
  assign Product1_4_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1207:1204]));
  assign Product1_5_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1463:1460]));
  assign Product1_6_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1719:1716]));
  assign Product1_7_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[2999:2996]));
  assign Product1_12_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3255:3252]));
  assign Product1_13_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3511:3508]));
  assign Product1_14_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3767:3764]));
  assign Product1_15_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1975:1972]));
  assign Product1_8_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2231:2228]));
  assign Product1_9_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2487:2484]));
  assign Product1_10_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2743:2740]));
  assign Product1_11_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1 = Accum2_acc_661_nl + Product1_1_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_46_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 = (Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4027:4024]));
  assign Product1_16_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_676_nl = Product1_16_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[187:184]);
  assign Accum2_acc_676_nl = nl_Accum2_acc_676_nl[7:0];
  assign nl_Product1_1_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[187:184]));
  assign Product1_1_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[443:440]));
  assign Product1_2_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[699:696]));
  assign Product1_3_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[955:952]));
  assign Product1_4_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1211:1208]));
  assign Product1_5_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1467:1464]));
  assign Product1_6_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1723:1720]));
  assign Product1_7_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3003:3000]));
  assign Product1_12_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3259:3256]));
  assign Product1_13_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3515:3512]));
  assign Product1_14_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3771:3768]));
  assign Product1_15_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1979:1976]));
  assign Product1_8_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2235:2232]));
  assign Product1_9_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2491:2488]));
  assign Product1_10_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2747:2744]));
  assign Product1_11_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1 = Accum2_acc_676_nl + Product1_1_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_47_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 = (Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4031:4028]));
  assign Product1_16_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_691_nl = Product1_16_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[191:188]);
  assign Accum2_acc_691_nl = nl_Accum2_acc_691_nl[7:0];
  assign nl_Product1_1_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[191:188]));
  assign Product1_1_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[447:444]));
  assign Product1_2_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[703:700]));
  assign Product1_3_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[959:956]));
  assign Product1_4_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1215:1212]));
  assign Product1_5_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1471:1468]));
  assign Product1_6_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1727:1724]));
  assign Product1_7_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3007:3004]));
  assign Product1_12_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3263:3260]));
  assign Product1_13_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3519:3516]));
  assign Product1_14_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3775:3772]));
  assign Product1_15_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1983:1980]));
  assign Product1_8_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2239:2236]));
  assign Product1_9_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2495:2492]));
  assign Product1_10_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2751:2748]));
  assign Product1_11_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1 = Accum2_acc_691_nl + Product1_1_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_48_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 = (Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4035:4032]));
  assign Product1_16_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_706_nl = Product1_16_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[195:192]);
  assign Accum2_acc_706_nl = nl_Accum2_acc_706_nl[7:0];
  assign nl_Product1_1_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[195:192]));
  assign Product1_1_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[451:448]));
  assign Product1_2_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[707:704]));
  assign Product1_3_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[963:960]));
  assign Product1_4_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1219:1216]));
  assign Product1_5_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1475:1472]));
  assign Product1_6_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1731:1728]));
  assign Product1_7_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3011:3008]));
  assign Product1_12_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3267:3264]));
  assign Product1_13_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3523:3520]));
  assign Product1_14_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3779:3776]));
  assign Product1_15_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1987:1984]));
  assign Product1_8_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2243:2240]));
  assign Product1_9_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2499:2496]));
  assign Product1_10_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2755:2752]));
  assign Product1_11_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1 = Accum2_acc_706_nl + Product1_1_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_49_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 = (Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4039:4036]));
  assign Product1_16_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_721_nl = Product1_16_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[199:196]);
  assign Accum2_acc_721_nl = nl_Accum2_acc_721_nl[7:0];
  assign nl_Product1_1_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[199:196]));
  assign Product1_1_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[455:452]));
  assign Product1_2_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[711:708]));
  assign Product1_3_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[967:964]));
  assign Product1_4_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1223:1220]));
  assign Product1_5_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1479:1476]));
  assign Product1_6_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1735:1732]));
  assign Product1_7_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3015:3012]));
  assign Product1_12_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3271:3268]));
  assign Product1_13_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3527:3524]));
  assign Product1_14_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3783:3780]));
  assign Product1_15_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1991:1988]));
  assign Product1_8_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2247:2244]));
  assign Product1_9_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2503:2500]));
  assign Product1_10_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2759:2756]));
  assign Product1_11_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1 = Accum2_acc_721_nl + Product1_1_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_50_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 = (Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4043:4040]));
  assign Product1_16_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_736_nl = Product1_16_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[203:200]);
  assign Accum2_acc_736_nl = nl_Accum2_acc_736_nl[7:0];
  assign nl_Product1_1_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[203:200]));
  assign Product1_1_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[459:456]));
  assign Product1_2_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[715:712]));
  assign Product1_3_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[971:968]));
  assign Product1_4_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1227:1224]));
  assign Product1_5_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1483:1480]));
  assign Product1_6_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1739:1736]));
  assign Product1_7_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3019:3016]));
  assign Product1_12_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3275:3272]));
  assign Product1_13_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3531:3528]));
  assign Product1_14_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3787:3784]));
  assign Product1_15_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1995:1992]));
  assign Product1_8_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2251:2248]));
  assign Product1_9_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2507:2504]));
  assign Product1_10_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2763:2760]));
  assign Product1_11_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1 = Accum2_acc_736_nl + Product1_1_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_51_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 = (Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4047:4044]));
  assign Product1_16_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_751_nl = Product1_16_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[207:204]);
  assign Accum2_acc_751_nl = nl_Accum2_acc_751_nl[7:0];
  assign nl_Product1_1_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[207:204]));
  assign Product1_1_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[463:460]));
  assign Product1_2_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[719:716]));
  assign Product1_3_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[975:972]));
  assign Product1_4_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1231:1228]));
  assign Product1_5_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1487:1484]));
  assign Product1_6_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1743:1740]));
  assign Product1_7_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3023:3020]));
  assign Product1_12_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3279:3276]));
  assign Product1_13_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3535:3532]));
  assign Product1_14_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3791:3788]));
  assign Product1_15_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[1999:1996]));
  assign Product1_8_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2255:2252]));
  assign Product1_9_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2511:2508]));
  assign Product1_10_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2767:2764]));
  assign Product1_11_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1 = Accum2_acc_751_nl + Product1_1_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_52_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 = (Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4051:4048]));
  assign Product1_16_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_766_nl = Product1_16_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[211:208]);
  assign Accum2_acc_766_nl = nl_Accum2_acc_766_nl[7:0];
  assign nl_Product1_1_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[211:208]));
  assign Product1_1_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[467:464]));
  assign Product1_2_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[723:720]));
  assign Product1_3_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[979:976]));
  assign Product1_4_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1235:1232]));
  assign Product1_5_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1491:1488]));
  assign Product1_6_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1747:1744]));
  assign Product1_7_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3027:3024]));
  assign Product1_12_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3283:3280]));
  assign Product1_13_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3539:3536]));
  assign Product1_14_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3795:3792]));
  assign Product1_15_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2003:2000]));
  assign Product1_8_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2259:2256]));
  assign Product1_9_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2515:2512]));
  assign Product1_10_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2771:2768]));
  assign Product1_11_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1 = Accum2_acc_766_nl + Product1_1_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_53_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 = (Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4055:4052]));
  assign Product1_16_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_781_nl = Product1_16_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[215:212]);
  assign Accum2_acc_781_nl = nl_Accum2_acc_781_nl[7:0];
  assign nl_Product1_1_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[215:212]));
  assign Product1_1_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[471:468]));
  assign Product1_2_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[727:724]));
  assign Product1_3_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[983:980]));
  assign Product1_4_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1239:1236]));
  assign Product1_5_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1495:1492]));
  assign Product1_6_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1751:1748]));
  assign Product1_7_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3031:3028]));
  assign Product1_12_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3287:3284]));
  assign Product1_13_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3543:3540]));
  assign Product1_14_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3799:3796]));
  assign Product1_15_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2007:2004]));
  assign Product1_8_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2263:2260]));
  assign Product1_9_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2519:2516]));
  assign Product1_10_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2775:2772]));
  assign Product1_11_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1 = Accum2_acc_781_nl + Product1_1_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_54_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 = (Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4059:4056]));
  assign Product1_16_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_796_nl = Product1_16_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[219:216]);
  assign Accum2_acc_796_nl = nl_Accum2_acc_796_nl[7:0];
  assign nl_Product1_1_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[219:216]));
  assign Product1_1_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[475:472]));
  assign Product1_2_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[731:728]));
  assign Product1_3_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[987:984]));
  assign Product1_4_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1243:1240]));
  assign Product1_5_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1499:1496]));
  assign Product1_6_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1755:1752]));
  assign Product1_7_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3035:3032]));
  assign Product1_12_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3291:3288]));
  assign Product1_13_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3547:3544]));
  assign Product1_14_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3803:3800]));
  assign Product1_15_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2011:2008]));
  assign Product1_8_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2267:2264]));
  assign Product1_9_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2523:2520]));
  assign Product1_10_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2779:2776]));
  assign Product1_11_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1 = Accum2_acc_796_nl + Product1_1_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_55_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 = (Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4063:4060]));
  assign Product1_16_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_811_nl = Product1_16_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[223:220]);
  assign Accum2_acc_811_nl = nl_Accum2_acc_811_nl[7:0];
  assign nl_Product1_1_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[223:220]));
  assign Product1_1_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[479:476]));
  assign Product1_2_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[735:732]));
  assign Product1_3_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[991:988]));
  assign Product1_4_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1247:1244]));
  assign Product1_5_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1503:1500]));
  assign Product1_6_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1759:1756]));
  assign Product1_7_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3039:3036]));
  assign Product1_12_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3295:3292]));
  assign Product1_13_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3551:3548]));
  assign Product1_14_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3807:3804]));
  assign Product1_15_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2015:2012]));
  assign Product1_8_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2271:2268]));
  assign Product1_9_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2527:2524]));
  assign Product1_10_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2783:2780]));
  assign Product1_11_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1 = Accum2_acc_811_nl + Product1_1_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_56_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 = (Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4067:4064]));
  assign Product1_16_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_826_nl = Product1_16_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[227:224]);
  assign Accum2_acc_826_nl = nl_Accum2_acc_826_nl[7:0];
  assign nl_Product1_1_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[227:224]));
  assign Product1_1_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[483:480]));
  assign Product1_2_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[739:736]));
  assign Product1_3_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[995:992]));
  assign Product1_4_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1251:1248]));
  assign Product1_5_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1507:1504]));
  assign Product1_6_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1763:1760]));
  assign Product1_7_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3043:3040]));
  assign Product1_12_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3299:3296]));
  assign Product1_13_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3555:3552]));
  assign Product1_14_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3811:3808]));
  assign Product1_15_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2019:2016]));
  assign Product1_8_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2275:2272]));
  assign Product1_9_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2531:2528]));
  assign Product1_10_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2787:2784]));
  assign Product1_11_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1 = Accum2_acc_826_nl + Product1_1_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_57_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1 = (Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4071:4068]));
  assign Product1_16_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_841_nl = Product1_16_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[231:228]);
  assign Accum2_acc_841_nl = nl_Accum2_acc_841_nl[7:0];
  assign nl_Product1_1_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[231:228]));
  assign Product1_1_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[487:484]));
  assign Product1_2_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[743:740]));
  assign Product1_3_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[999:996]));
  assign Product1_4_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1255:1252]));
  assign Product1_5_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1511:1508]));
  assign Product1_6_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1767:1764]));
  assign Product1_7_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3047:3044]));
  assign Product1_12_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3303:3300]));
  assign Product1_13_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3559:3556]));
  assign Product1_14_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3815:3812]));
  assign Product1_15_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2023:2020]));
  assign Product1_8_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2279:2276]));
  assign Product1_9_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2535:2532]));
  assign Product1_10_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2791:2788]));
  assign Product1_11_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1 = Accum2_acc_841_nl + Product1_1_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_58_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1 = (Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4075:4072]));
  assign Product1_16_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_856_nl = Product1_16_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[235:232]);
  assign Accum2_acc_856_nl = nl_Accum2_acc_856_nl[7:0];
  assign nl_Product1_1_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[235:232]));
  assign Product1_1_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[491:488]));
  assign Product1_2_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[747:744]));
  assign Product1_3_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1003:1000]));
  assign Product1_4_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1259:1256]));
  assign Product1_5_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1515:1512]));
  assign Product1_6_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1771:1768]));
  assign Product1_7_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3051:3048]));
  assign Product1_12_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3307:3304]));
  assign Product1_13_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3563:3560]));
  assign Product1_14_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3819:3816]));
  assign Product1_15_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2027:2024]));
  assign Product1_8_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2283:2280]));
  assign Product1_9_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2539:2536]));
  assign Product1_10_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2795:2792]));
  assign Product1_11_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1 = Accum2_acc_856_nl + Product1_1_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_59_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1 = (Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4079:4076]));
  assign Product1_16_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_871_nl = Product1_16_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[239:236]);
  assign Accum2_acc_871_nl = nl_Accum2_acc_871_nl[7:0];
  assign nl_Product1_1_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[239:236]));
  assign Product1_1_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[495:492]));
  assign Product1_2_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[751:748]));
  assign Product1_3_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1007:1004]));
  assign Product1_4_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1263:1260]));
  assign Product1_5_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1519:1516]));
  assign Product1_6_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1775:1772]));
  assign Product1_7_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3055:3052]));
  assign Product1_12_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3311:3308]));
  assign Product1_13_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3567:3564]));
  assign Product1_14_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3823:3820]));
  assign Product1_15_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2031:2028]));
  assign Product1_8_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2287:2284]));
  assign Product1_9_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2543:2540]));
  assign Product1_10_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2799:2796]));
  assign Product1_11_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1 = Accum2_acc_871_nl + Product1_1_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_60_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1 = (Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4083:4080]));
  assign Product1_16_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_886_nl = Product1_16_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[243:240]);
  assign Accum2_acc_886_nl = nl_Accum2_acc_886_nl[7:0];
  assign nl_Product1_1_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[243:240]));
  assign Product1_1_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[499:496]));
  assign Product1_2_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[755:752]));
  assign Product1_3_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1011:1008]));
  assign Product1_4_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1267:1264]));
  assign Product1_5_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1523:1520]));
  assign Product1_6_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1779:1776]));
  assign Product1_7_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3059:3056]));
  assign Product1_12_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3315:3312]));
  assign Product1_13_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3571:3568]));
  assign Product1_14_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3827:3824]));
  assign Product1_15_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2035:2032]));
  assign Product1_8_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2291:2288]));
  assign Product1_9_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2547:2544]));
  assign Product1_10_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2803:2800]));
  assign Product1_11_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1 = Accum2_acc_886_nl + Product1_1_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_61_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1 = (Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4087:4084]));
  assign Product1_16_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_901_nl = Product1_16_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[247:244]);
  assign Accum2_acc_901_nl = nl_Accum2_acc_901_nl[7:0];
  assign nl_Product1_1_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[247:244]));
  assign Product1_1_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[503:500]));
  assign Product1_2_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[759:756]));
  assign Product1_3_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1015:1012]));
  assign Product1_4_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1271:1268]));
  assign Product1_5_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1527:1524]));
  assign Product1_6_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1783:1780]));
  assign Product1_7_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3063:3060]));
  assign Product1_12_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3319:3316]));
  assign Product1_13_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3575:3572]));
  assign Product1_14_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3831:3828]));
  assign Product1_15_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2039:2036]));
  assign Product1_8_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2295:2292]));
  assign Product1_9_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2551:2548]));
  assign Product1_10_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2807:2804]));
  assign Product1_11_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1 = Accum2_acc_901_nl + Product1_1_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_62_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1 = (Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4091:4088]));
  assign Product1_16_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_916_nl = Product1_16_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[251:248]);
  assign Accum2_acc_916_nl = nl_Accum2_acc_916_nl[7:0];
  assign nl_Product1_1_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[251:248]));
  assign Product1_1_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[507:504]));
  assign Product1_2_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[763:760]));
  assign Product1_3_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1019:1016]));
  assign Product1_4_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1275:1272]));
  assign Product1_5_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1531:1528]));
  assign Product1_6_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1787:1784]));
  assign Product1_7_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3067:3064]));
  assign Product1_12_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3323:3320]));
  assign Product1_13_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3579:3576]));
  assign Product1_14_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3835:3832]));
  assign Product1_15_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2043:2040]));
  assign Product1_8_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2299:2296]));
  assign Product1_9_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2555:2552]));
  assign Product1_10_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2811:2808]));
  assign Product1_11_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1 = Accum2_acc_916_nl + Product1_1_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_63_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 = (Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1[6:3]!=4'b0000);
  assign nl_Product1_16_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4095:4092]));
  assign Product1_16_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum2_acc_931_nl = Product1_16_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_4_8(b2_rsci_idat[255:252]);
  assign Accum2_acc_931_nl = nl_Accum2_acc_931_nl[7:0];
  assign nl_Product1_1_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[255:252]));
  assign Product1_1_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_2_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[511:508]));
  assign Product1_2_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_3_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[767:764]));
  assign Product1_3_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_4_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1023:1020]));
  assign Product1_4_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_5_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1279:1276]));
  assign Product1_5_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_6_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1535:1532]));
  assign Product1_6_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_7_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1791:1788]));
  assign Product1_7_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_12_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3071:3068]));
  assign Product1_12_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_13_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3327:3324]));
  assign Product1_13_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_14_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3583:3580]));
  assign Product1_14_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_15_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[3839:3836]));
  assign Product1_15_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_8_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2047:2044]));
  assign Product1_8_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_9_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2303:2300]));
  assign Product1_9_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_10_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2559:2556]));
  assign Product1_10_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Product1_11_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2815:2812]));
  assign Product1_11_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[7:0];
  assign nl_Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1 = Accum2_acc_931_nl + Product1_1_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_4_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_6_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_7_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_12_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_13_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_64_operator_4_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1 = nl_Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1[7:0];
  assign nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[739:736]));
  assign Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[703:700]));
  assign Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[643:640]));
  assign Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[607:604]));
  assign Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[691:688]));
  assign Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[655:652]));
  assign Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[67:64]));
  assign Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[79:76]));
  assign Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[19:16]));
  assign Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[31:28]));
  assign Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[43:40]));
  assign Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[55:52]));
  assign Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[595:592]));
  assign Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[559:556]));
  assign Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[571:568]));
  assign Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[535:532]));
  assign Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum2_1_acc_192_nl = conv_s2s_4_5(b5_rsci_idat[7:4]) + conv_s2s_4_5(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1[4:1]);
  assign Accum2_1_acc_192_nl = nl_Accum2_1_acc_192_nl[4:0];
  assign nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[547:544]));
  assign Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[523:520]));
  assign Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[751:748]));
  assign Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[499:496]));
  assign Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[511:508]));
  assign Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[763:760]));
  assign Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[727:724]));
  assign Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[715:712]));
  assign Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[679:676]));
  assign Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[667:664]));
  assign Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[631:628]));
  assign Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[619:616]));
  assign Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[583:580]));
  assign Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[91:88]));
  assign Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[103:100]));
  assign Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum2_1_acc_127_nl = conv_s2s_5_10(readslicef_12_5_7(Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_6_10({Accum2_1_acc_192_nl , (Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1[0])})
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum2_1_acc_127_nl = nl_Accum2_1_acc_127_nl[9:0];
  assign nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[259:256]));
  assign Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[271:268]));
  assign Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[211:208]));
  assign Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[223:220]));
  assign Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[115:112]));
  assign Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[127:124]));
  assign Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[139:136]));
  assign Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[151:148]));
  assign Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[163:160]));
  assign Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[175:172]));
  assign Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[187:184]));
  assign Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[199:196]));
  assign Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[307:304]));
  assign Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[319:316]));
  assign Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[331:328]));
  assign Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[343:340]));
  assign Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[355:352]));
  assign Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[367:364]));
  assign Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[379:376]));
  assign Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[391:388]));
  assign Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[451:448]));
  assign Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[463:460]));
  assign Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[475:472]));
  assign Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[487:484]));
  assign Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[403:400]));
  assign Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[415:412]));
  assign Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[427:424]));
  assign Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[439:436]));
  assign Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[235:232]));
  assign Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[247:244]));
  assign Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[283:280]));
  assign Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[295:292]));
  assign Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1 = Accum2_1_acc_127_nl
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1 = nl_Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1[9:0];
  assign nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[719:716]));
  assign Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[731:728]));
  assign Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[623:620]));
  assign Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[635:632]));
  assign Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[671:668]));
  assign Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[683:680]));
  assign Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[59:56]));
  assign Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[71:68]));
  assign Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({layer4_out_conc_4_7 , layer4_out_conc_4_6_5 , ({{3{layer4_out_0_1_lpi_1_dfm_1}},
      layer4_out_0_1_lpi_1_dfm_1}) , layer4_out_0_1_lpi_1_dfm_1})) * $signed((w5_rsci_idat[11:8]));
  assign Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[23:20]));
  assign Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[35:32]));
  assign Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[47:44]));
  assign Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[575:572]));
  assign Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[587:584]));
  assign Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[551:548]));
  assign Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[563:560]));
  assign Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum2_1_acc_193_nl = conv_s2s_4_5(Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1[4:1])
      + conv_s2s_4_5(b5_rsci_idat[11:8]);
  assign Accum2_1_acc_193_nl = nl_Accum2_1_acc_193_nl[4:0];
  assign nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[527:524]));
  assign Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[539:536]));
  assign Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[743:740]));
  assign Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[491:488]));
  assign Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[503:500]));
  assign Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[755:752]));
  assign Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[767:764]));
  assign Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[695:692]));
  assign Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[707:704]));
  assign Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[647:644]));
  assign Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[659:656]));
  assign Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[599:596]));
  assign Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[611:608]));
  assign Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[83:80]));
  assign Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[95:92]));
  assign Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum2_1_acc_190_nl = conv_s2s_5_10(readslicef_12_5_7(Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_6_10({Accum2_1_acc_193_nl , (Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1[0])})
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum2_1_acc_190_nl = nl_Accum2_1_acc_190_nl[9:0];
  assign nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[251:248]));
  assign Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[263:260]));
  assign Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[203:200]));
  assign Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[215:212]));
  assign Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[107:104]));
  assign Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[119:116]));
  assign Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[131:128]));
  assign Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[143:140]));
  assign Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[155:152]));
  assign Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[167:164]));
  assign Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[179:176]));
  assign Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[191:188]));
  assign Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[299:296]));
  assign Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[311:308]));
  assign Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[323:320]));
  assign Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[335:332]));
  assign Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[347:344]));
  assign Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[359:356]));
  assign Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[371:368]));
  assign Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[383:380]));
  assign Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[443:440]));
  assign Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[455:452]));
  assign Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[467:464]));
  assign Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[479:476]));
  assign Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[395:392]));
  assign Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[407:404]));
  assign Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[419:416]));
  assign Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[431:428]));
  assign Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[227:224]));
  assign Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[239:236]));
  assign Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[275:272]));
  assign Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[287:284]));
  assign Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1 = Accum2_1_acc_190_nl
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1 = nl_Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1[9:0];
  assign nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[735:732]));
  assign Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[699:696]));
  assign Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[639:636]));
  assign Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[603:600]));
  assign Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[687:684]));
  assign Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[651:648]));
  assign Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[63:60]));
  assign Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[75:72]));
  assign Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[15:12]));
  assign Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[27:24]));
  assign Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[39:36]));
  assign Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[51:48]));
  assign Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[591:588]));
  assign Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[555:552]));
  assign Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[567:564]));
  assign Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[531:528]));
  assign Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum2_1_acc_191_nl = conv_s2s_4_5(b5_rsci_idat[3:0]) + conv_s2s_4_5(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1[4:1]);
  assign Accum2_1_acc_191_nl = nl_Accum2_1_acc_191_nl[4:0];
  assign nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[543:540]));
  assign Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[519:516]));
  assign Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[747:744]));
  assign Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[495:492]));
  assign Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[507:504]));
  assign Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[759:756]));
  assign Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[723:720]));
  assign Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[711:708]));
  assign Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[675:672]));
  assign Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[663:660]));
  assign Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[627:624]));
  assign Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[615:612]));
  assign Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[579:576]));
  assign Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[87:84]));
  assign Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[99:96]));
  assign Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum2_1_acc_nl = conv_s2s_5_10(readslicef_12_5_7(Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_6_10({Accum2_1_acc_191_nl , (Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1[0])})
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum2_1_acc_nl = nl_Accum2_1_acc_nl[9:0];
  assign nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[255:252]));
  assign Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[267:264]));
  assign Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[207:204]));
  assign Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[219:216]));
  assign Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[111:108]));
  assign Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[123:120]));
  assign Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[135:132]));
  assign Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[147:144]));
  assign Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[159:156]));
  assign Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[171:168]));
  assign Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[183:180]));
  assign Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[195:192]));
  assign Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[303:300]));
  assign Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[315:312]));
  assign Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[327:324]));
  assign Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[339:336]));
  assign Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[351:348]));
  assign Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[363:360]));
  assign Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[375:372]));
  assign Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[387:384]));
  assign Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[447:444]));
  assign Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[459:456]));
  assign Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[471:468]));
  assign Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[483:480]));
  assign Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[399:396]));
  assign Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[411:408]));
  assign Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[423:420]));
  assign Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[435:432]));
  assign Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[231:228]));
  assign Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[243:240]));
  assign Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[279:276]));
  assign Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[291:288]));
  assign Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign nl_Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1 = Accum2_1_acc_nl +
      conv_s2s_5_10(readslicef_12_5_7(Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_5_10(readslicef_12_5_7(Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1 = nl_Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1[9:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_8_1;
  assign nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_7
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_6_5 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[515:512]));
  assign Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1
      = readslicef_12_5_7(Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign layer4_out_0_1_lpi_1_dfm_1 = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1
      & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_8_1;
  assign nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({layer4_out_conc_4_7 , layer4_out_conc_4_6_5 , ({{3{layer4_out_0_1_lpi_1_dfm_1}},
      layer4_out_0_1_lpi_1_dfm_1}) , layer4_out_0_1_lpi_1_dfm_1})) * $signed((w5_rsci_idat[7:4]));
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1
      = readslicef_12_5_7(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_8_9({layer4_out_conc_4_7 , layer4_out_conc_4_6_5 , ({{3{layer4_out_0_1_lpi_1_dfm_1}},
      layer4_out_0_1_lpi_1_dfm_1}) , layer4_out_0_1_lpi_1_dfm_1})) * $signed((w5_rsci_idat[3:0]));
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[11:0];
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_11_7_1
      = readslicef_12_5_7(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl =  -conv_s2s_8_9(Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl =  -conv_s2s_8_9(Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl =  -conv_s2s_8_9(Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl =  -conv_s2s_8_9(Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl =  -conv_s2s_8_9(Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl =  -conv_s2s_8_9(Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl =  -conv_s2s_8_9(Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl =  -conv_s2s_8_9(Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl =  -conv_s2s_8_9(Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl =  -conv_s2s_8_9(Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl =  -conv_s2s_8_9(Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl =  -conv_s2s_8_9(Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl =  -conv_s2s_8_9(Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl =  -conv_s2s_8_9(Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl =  -conv_s2s_8_9(Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl =  -conv_s2s_8_9(Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl =  -conv_s2s_8_9(Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl =  -conv_s2s_8_9(Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl =  -conv_s2s_8_9(Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl =  -conv_s2s_8_9(Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl =  -conv_s2s_8_9(Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl =  -conv_s2s_8_9(Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl =  -conv_s2s_8_9(Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl =  -conv_s2s_8_9(Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl =  -conv_s2s_8_9(Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl =  -conv_s2s_8_9(Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl =  -conv_s2s_8_9(Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl =  -conv_s2s_8_9(Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl =  -conv_s2s_8_9(Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl =  -conv_s2s_8_9(Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl =  -conv_s2s_8_9(Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl =  -conv_s2s_8_9(Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl =  -conv_s2s_8_9(Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl =  -conv_s2s_8_9(Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl =  -conv_s2s_8_9(Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl =  -conv_s2s_8_9(Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl =  -conv_s2s_8_9(Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl =  -conv_s2s_8_9(Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl =  -conv_s2s_8_9(Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl =  -conv_s2s_8_9(Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl =  -conv_s2s_8_9(Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl =  -conv_s2s_8_9(Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl =  -conv_s2s_8_9(Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl =  -conv_s2s_8_9(Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl =  -conv_s2s_8_9(Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl =  -conv_s2s_8_9(Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl =  -conv_s2s_8_9(Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl =  -conv_s2s_8_9(Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl =  -conv_s2s_8_9(Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl =  -conv_s2s_8_9(Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl =  -conv_s2s_8_9(Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl =  -conv_s2s_8_9(Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl =  -conv_s2s_8_9(Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl =  -conv_s2s_8_9(Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl =  -conv_s2s_8_9(Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl =  -conv_s2s_8_9(Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl =  -conv_s2s_8_9(Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl =  -conv_s2s_8_9(Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl =  -conv_s2s_8_9(Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl =  -conv_s2s_8_9(Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl =  -conv_s2s_8_9(Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl =  -conv_s2s_8_9(Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl =  -conv_s2s_8_9(Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl =  -conv_s2s_8_9(Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl[8:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_8_1 = readslicef_9_1_8(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_7 = ((Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_41_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_192_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_7 = ((Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_42_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_194_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_7 = ((Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_62_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_196_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_7 = ((Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_63_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_198_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_7 = ((Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_64_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_200_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_7 = ((Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_60_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_202_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_7 = ((Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_61_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_7 = ((Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_58_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_7 = ((Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_59_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_7 = ((Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_56_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_7 = ((Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_57_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_7 = ((Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_54_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_7 = ((Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_55_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_7 = ((Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_52_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_7 = ((Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_53_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_7 = ((Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_50_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_7 = ((Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_51_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_7 = ((Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_48_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_7 = ((Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_49_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_7 = ((Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_46_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_7 = ((Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_47_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_7 = ((Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_44_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_7 = ((Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_45_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_8_1);
  assign layer4_out_conc_4_7 = ((Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1[2]) |
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_1_Accum2_acc_1_psp_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1);
  assign layer4_out_conc_4_6_5 = MUX_v_2_2_2(2'b00, nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_7 = ((Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_2_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_7 = ((Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_3_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_7 = ((Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_4_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_7 = ((Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_5_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_7 = ((Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_6_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_7 = ((Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_7_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_7 = ((Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_8_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_7 = ((Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_9_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_7 = ((Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_10_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_7 = ((Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_11_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_7 = ((Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_12_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_7 = ((Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_13_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_7 = ((Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_14_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_7 = ((Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_15_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_7 = ((Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_16_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_7 = ((Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_17_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_7 = ((Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_18_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_7 = ((Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_19_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_7 = ((Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_20_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_7 = ((Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_21_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_7 = ((Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_22_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_7 = ((Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_23_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_7 = ((Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_24_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_7 = ((Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_25_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_7 = ((Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_26_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_7 = ((Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_27_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_7 = ((Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_28_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_7 = ((Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_29_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_7 = ((Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_30_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_7 = ((Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_31_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_7 = ((Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_32_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_7 = ((Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_33_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_7 = ((Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_34_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_7 = ((Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_35_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_7 = ((Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_36_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_7 = ((Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_37_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_7 = ((Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_38_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_7 = ((Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_39_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_7 = ((Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_40_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_8_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_7 = ((Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1[2])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_8_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl
      = MUX_v_2_2_2((Accum1_16_Accum2_43_Accum2_acc_1_ncse_sva_1[1:0]), 2'b11, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_6_5 = MUX_v_2_2_2(2'b00,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_3_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_8_1);
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat <= 2'b00;
    end
    else begin
      layer7_out_rsci_idat <= ~(MUX_v_2_2_2(argmax_else_mux_nl, 2'b11, argmax_if_argmax_if_argmax_if_nor_nl));
    end
  end
  assign nl_argmax_else_aelse_acc_nl = conv_s2u_10_11(Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1)
      - conv_s2u_10_11(Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1);
  assign argmax_else_aelse_acc_nl = nl_argmax_else_aelse_acc_nl[10:0];
  assign nl_argmax_else_if_acc_nl = conv_s2u_10_11(Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1)
      - conv_s2u_10_11(Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1);
  assign argmax_else_if_acc_nl = nl_argmax_else_if_acc_nl[10:0];
  assign argmax_else_if_argmax_else_if_argmax_else_if_nor_nl = ~((readslicef_11_1_10(argmax_else_aelse_acc_nl))
      | (readslicef_11_1_10(argmax_else_if_acc_nl)));
  assign argmax_else_mux_nl = MUX_v_2_2_2(2'b01, 2'b10, argmax_else_if_argmax_else_if_argmax_else_if_nor_nl);
  assign nl_argmax_aelse_acc_nl = conv_s2u_10_11(Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1)
      - conv_s2u_10_11(Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1);
  assign argmax_aelse_acc_nl = nl_argmax_aelse_acc_nl[10:0];
  assign nl_argmax_if_acc_nl = conv_s2u_10_11(Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1)
      - conv_s2u_10_11(Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1);
  assign argmax_if_acc_nl = nl_argmax_if_acc_nl[10:0];
  assign argmax_if_argmax_if_argmax_if_nor_nl = ~((readslicef_11_1_10(argmax_aelse_acc_nl))
      | (readslicef_11_1_10(argmax_if_acc_nl)));

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] readslicef_12_5_7;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_12_5_7 = tmp[4:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] conv_s2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2s_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [7:0] conv_s2s_4_8 ;
    input [3:0]  vector ;
  begin
    conv_s2s_4_8 = {{4{vector[3]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_5_10 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_10 = {{5{vector[4]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_6_10 ;
    input [5:0]  vector ;
  begin
    conv_s2s_6_10 = {{4{vector[5]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    myproject
// ------------------------------------------------------------------


module myproject (
  clk, rst, input_1_rsc_dat, layer7_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [95:0] input_1_rsc_dat;
  output [1:0] layer7_out_rsc_dat;
  input [4095:0] w2_rsc_dat;
  input [255:0] b2_rsc_dat;
  input [767:0] w5_rsc_dat;
  input [11:0] b5_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  converterBlock_myproject_core myproject_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .w2_rsc_dat(w2_rsc_dat),
      .b2_rsc_dat(b2_rsc_dat),
      .w5_rsc_dat(w5_rsc_dat),
      .b5_rsc_dat(b5_rsc_dat)
    );
endmodule



