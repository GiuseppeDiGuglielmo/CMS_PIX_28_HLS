
//------> ./myproject_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module converterBlock_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./myproject_ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module converterBlock_ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./myproject.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
// 
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Mon Oct 24 21:18:19 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core
// ------------------------------------------------------------------


module converterBlock_myproject_core (
  clk, rst, input_1_rsc_dat, layer6_out_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer6_out_rsc_dat;


  // Interconnect Declarations
  wire [223:0] input_1_rsci_idat;
  reg [15:0] layer6_out_rsci_idat_47_32;
  wire [18:0] nl_layer6_out_rsci_idat_47_32;
  reg [15:0] layer6_out_rsci_idat_31_16;
  wire [16:0] nl_layer6_out_rsci_idat_31_16;
  reg [14:0] layer6_out_rsci_idat_14_0;
  wire [16:0] nl_layer6_out_rsci_idat_14_0;
  wire [15:0] Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1;
  wire [15:0] Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1;
  wire [19:0] nl_Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1;
  wire [17:0] nl_Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1;
  wire [18:0] nl_Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1;
  wire [19:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1;
  wire [19:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1;
  wire [19:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1;
  wire [19:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1;
  wire [19:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1;
  wire [17:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1;
  wire [18:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [11:0] Product2_1_acc_722_cse_1;
  wire [12:0] nl_Product2_1_acc_722_cse_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire [8:0] layer4_out_0_9_1_lpi_1_dfm_1;
  wire layer4_out_0_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [7:0] nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1;
  wire [8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [8:0] nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1;
  wire [9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_9_lpi_1_dfm_1;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_8_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_0_lpi_1_dfm_1;
  wire [6:0] Accum2_acc_1558_cse_1;
  wire [7:0] nl_Accum2_acc_1558_cse_1;
  wire [15:0] Product2_acc_792_cse_sva_1;
  wire [16:0] nl_Product2_acc_792_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_532_cse_sva_1;
  wire [16:0] nl_Product2_acc_532_cse_sva_1;
  wire [13:0] Accum2_acc_1313_cse_1;
  wire [14:0] nl_Accum2_acc_1313_cse_1;
  wire [15:0] Accum2_acc_411_cse_1;
  wire [16:0] nl_Accum2_acc_411_cse_1;
  wire [15:0] Product2_acc_308_cse_sva_1;
  wire [16:0] nl_Product2_acc_308_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1;
  wire [15:0] Product2_acc_195_cse_sva_1;
  wire [16:0] nl_Product2_acc_195_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_124_cse_sva_1;
  wire [16:0] nl_Product2_acc_124_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_368_cse_sva_1;
  wire [16:0] nl_Product2_acc_368_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] Accum2_acc_1028_cse_1;
  wire [14:0] nl_Accum2_acc_1028_cse_1;
  wire [13:0] Accum2_acc_476_cse_1;
  wire [14:0] nl_Accum2_acc_476_cse_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_370_cse_sva_1;
  wire [16:0] nl_Product2_acc_370_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1;
  wire [15:0] Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Accum2_acc_1066_cse_1;
  wire [16:0] nl_Accum2_acc_1066_cse_1;
  wire [15:0] Product2_acc_797_cse_sva_1;
  wire [16:0] nl_Product2_acc_797_cse_sva_1;
  wire [15:0] Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_204_cse_sva_1;
  wire [16:0] nl_Product2_acc_204_cse_sva_1;
  wire [15:0] Product2_acc_943_cse_sva_1;
  wire [16:0] nl_Product2_acc_943_cse_sva_1;
  wire [15:0] Product2_acc_730_cse_sva_1;
  wire [16:0] nl_Product2_acc_730_cse_sva_1;
  wire [15:0] Product2_acc_667_cse_sva_1;
  wire [16:0] nl_Product2_acc_667_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1;
  wire [13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1;
  wire [15:0] Accum2_acc_399_cse_1;
  wire [16:0] nl_Accum2_acc_399_cse_1;
  wire [15:0] Product2_acc_867_cse_sva_1;
  wire [16:0] nl_Product2_acc_867_cse_sva_1;
  wire [12:0] Accum2_acc_1120_cse_1;
  wire [13:0] nl_Accum2_acc_1120_cse_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_609_cse_sva_1;
  wire [16:0] nl_Product2_acc_609_cse_sva_1;
  wire [15:0] Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] Accum2_acc_1027_cse_1;
  wire [14:0] nl_Accum2_acc_1027_cse_1;
  wire [12:0] Accum2_acc_825_cse_1;
  wire [13:0] nl_Accum2_acc_825_cse_1;
  wire [15:0] Product2_acc_127_cse_sva_1;
  wire [16:0] nl_Product2_acc_127_cse_sva_1;
  wire [15:0] Accum2_acc_426_cse_1;
  wire [16:0] nl_Accum2_acc_426_cse_1;
  wire [15:0] Product2_acc_214_cse_sva_1;
  wire [16:0] nl_Product2_acc_214_cse_sva_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] Accum2_acc_727_cse_1;
  wire [14:0] nl_Accum2_acc_727_cse_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_665_cse_sva_1;
  wire [16:0] nl_Product2_acc_665_cse_sva_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] Accum2_acc_992_cse_1;
  wire [14:0] nl_Accum2_acc_992_cse_1;
  wire [15:0] Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Accum2_acc_766_cse_1;
  wire [16:0] nl_Accum2_acc_766_cse_1;
  wire [13:0] Accum2_acc_295_cse_1;
  wire [14:0] nl_Accum2_acc_295_cse_1;
  wire [15:0] Product2_acc_970_cse_sva_1;
  wire [16:0] nl_Product2_acc_970_cse_sva_1;
  wire [14:0] Accum2_acc_447_cse_1;
  wire [15:0] nl_Accum2_acc_447_cse_1;
  wire [15:0] Product2_acc_538_cse_sva_1;
  wire [16:0] nl_Product2_acc_538_cse_sva_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [12:0] Accum2_acc_532_cse_1;
  wire [13:0] nl_Accum2_acc_532_cse_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_936_cse_sva_1;
  wire [16:0] nl_Product2_acc_936_cse_sva_1;
  wire [12:0] Accum2_acc_306_cse_1;
  wire [13:0] nl_Accum2_acc_306_cse_1;
  wire [13:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Accum2_acc_590_cse_1;
  wire [16:0] nl_Accum2_acc_590_cse_1;
  wire [13:0] Accum2_acc_534_cse_1;
  wire [14:0] nl_Accum2_acc_534_cse_1;
  wire [14:0] Accum2_acc_343_cse_1;
  wire [15:0] nl_Accum2_acc_343_cse_1;
  wire [15:0] Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [16:0] nl_Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_794_cse_sva_1;
  wire [16:0] nl_Product2_acc_794_cse_sva_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_382_cse_sva_1;
  wire [16:0] nl_Product2_acc_382_cse_sva_1;
  wire [13:0] Accum2_acc_635_cse_1;
  wire [14:0] nl_Accum2_acc_635_cse_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Product2_acc_743_cse_sva_1;
  wire [16:0] nl_Product2_acc_743_cse_sva_1;
  wire [14:0] Accum2_acc_457_cse_1;
  wire [15:0] nl_Accum2_acc_457_cse_1;
  wire [15:0] Product2_acc_459_cse_sva_1;
  wire [16:0] nl_Product2_acc_459_cse_sva_1;
  wire [14:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [13:0] Accum2_acc_387_cse_1;
  wire [14:0] nl_Accum2_acc_387_cse_1;
  wire [15:0] nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  wire [15:0] Accum2_acc_285_cse_1;
  wire [16:0] nl_Accum2_acc_285_cse_1;
  wire [15:0] Accum2_acc_261_cse_1;
  wire [16:0] nl_Accum2_acc_261_cse_1;
  wire [15:0] Accum2_acc_215_cse_1;
  wire [16:0] nl_Accum2_acc_215_cse_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_not_279;
  wire Product2_1_not_911;
  wire Product2_1_not_941;
  wire Product2_1_not_943;
  wire Product2_1_not_949;
  wire Product2_1_not_963;
  wire [15:0] Accum2_acc_1648;
  wire [16:0] nl_Accum2_acc_1648;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [8:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_0;
  wire [5:0] Accum2_Accum2_conc_111_12_7;
  wire [6:0] nl_Accum2_Accum2_conc_111_12_7;
  wire [3:0] Accum2_Accum2_conc_113_12_9;
  wire [4:0] nl_Accum2_Accum2_conc_113_12_9;
  wire [5:0] Accum2_Accum2_conc_115_12_7;
  wire [6:0] nl_Accum2_Accum2_conc_115_12_7;
  wire [6:0] Accum2_Accum2_conc_117_12_6;
  wire [7:0] nl_Accum2_Accum2_conc_117_12_6;
  wire [6:0] Accum2_Accum2_conc_119_12_6;
  wire [7:0] nl_Accum2_Accum2_conc_119_12_6;
  wire [4:0] Accum2_Accum2_conc_121_12_8;
  wire [5:0] nl_Accum2_Accum2_conc_121_12_8;
  wire [5:0] Accum2_Accum2_conc_123_12_7;
  wire [6:0] nl_Accum2_Accum2_conc_123_12_7;
  wire [6:0] Accum2_Accum2_conc_125_12_6;
  wire [7:0] nl_Accum2_Accum2_conc_125_12_6;
  wire [5:0] Accum2_Accum2_conc_127_12_7;
  wire [6:0] nl_Accum2_Accum2_conc_127_12_7;
  wire [4:0] Accum2_Accum2_conc_129_12_8;
  wire [5:0] nl_Accum2_Accum2_conc_129_12_8;
  wire [10:0] Product2_1_acc_415_itm_13_3_1;
  wire [10:0] Product2_1_acc_418_itm_12_2_1;
  wire [10:0] Product2_1_acc_423_itm_12_2_1;
  wire [10:0] Product2_1_acc_424_itm_13_3_1;
  wire [10:0] Product2_1_acc_425_itm_13_3_1;
  wire [10:0] Product2_1_acc_428_itm_12_2_1;
  wire [10:0] Product2_1_acc_429_itm_12_2_1;
  wire [10:0] Product2_1_acc_430_itm_13_3_1;
  wire [10:0] Product2_1_acc_431_itm_12_2_1;
  wire [7:0] Product2_1_acc_67_itm_11_4_1;
  wire [9:0] Product2_1_acc_384_itm_10_1_1;
  wire [10:0] Product2_1_acc_396_itm_12_2_1;
  wire [7:0] Product2_1_acc_76_itm_11_4_1;
  wire [10:0] Product2_1_acc_391_itm_12_2_1;
  wire [10:0] Product2_1_acc_393_itm_12_2_1;
  wire [10:0] Product2_1_acc_399_itm_12_2_1;
  wire [8:0] Product2_1_acc_478_itm_10_2_1;
  wire [8:0] Product2_1_acc_72_itm_11_3_1;
  wire [7:0] Product2_1_acc_241_itm_11_4_1;
  wire [9:0] Product2_1_acc_469_itm_10_1_1;
  wire [9:0] Product2_1_acc_8_itm_11_2_1;
  wire [10:0] Product2_1_acc_410_itm_13_3_1;
  wire [10:0] Product2_1_acc_411_itm_13_3_1;
  wire [10:0] Product2_1_acc_414_itm_12_2_1;
  wire [10:0] Product2_1_acc_644_itm_13_3_1;
  wire [10:0] Product2_1_acc_645_itm_12_2_1;
  wire [10:0] Product2_1_acc_633_itm_12_2_1;
  wire [10:0] Product2_1_acc_634_itm_12_2_1;
  wire [10:0] Product2_1_acc_636_itm_12_2_1;
  wire [10:0] Product2_1_acc_638_itm_12_2_1;
  wire [10:0] Product2_1_acc_641_itm_12_2_1;
  wire [10:0] Product2_1_acc_642_itm_12_2_1;
  wire [7:0] Product2_1_acc_79_itm_11_4_1;
  wire [10:0] Product2_1_acc_643_itm_13_3_1;
  wire [10:0] Product2_1_acc_476_itm_13_3_1;
  wire [10:0] Product2_1_acc_477_itm_13_3_1;
  wire [10:0] Product2_1_acc_480_itm_13_3_1;
  wire [10:0] Product2_1_acc_483_itm_13_3_1;
  wire [10:0] Product2_1_acc_484_itm_12_2_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire [10:0] Product2_1_acc_450_itm_12_2_1;
  wire [10:0] Product2_1_acc_462_itm_12_2_1;
  wire [10:0] Product2_1_acc_464_itm_12_2_1;
  wire [10:0] Product2_1_acc_454_itm_12_2_1;
  wire [10:0] Product2_1_acc_455_itm_12_2_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire [10:0] Product2_1_acc_466_itm_13_3_1;
  wire [10:0] Product2_1_acc_467_itm_12_2_1;
  wire [10:0] Product2_1_acc_468_itm_13_3_1;
  wire [10:0] Product2_1_acc_473_itm_13_3_1;
  wire [10:0] Product2_1_acc_474_itm_13_3_1;
  wire [10:0] Product2_1_acc_475_itm_12_2_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire [14:0] Product2_acc_1027_itm_16_2_1;
  wire [15:0] Product2_acc_478_itm_17_2_1;
  wire [15:0] Product2_acc_377_itm_17_2_1;
  wire [15:0] Product2_acc_946_itm_18_3_1;
  wire [15:0] Product2_acc_1064_itm_16_1_1;
  wire [15:0] Product2_acc_1134_itm_16_1_1;
  wire [15:0] Product2_acc_1034_itm_16_1_1;
  wire [15:0] Product2_acc_297_itm_17_2_1;
  wire [15:0] Product2_acc_75_itm_19_4_1;
  wire [15:0] Product2_acc_728_itm_18_3_1;
  wire [15:0] Product2_acc_834_itm_19_4_1;
  wire [15:0] Product2_acc_934_itm_17_2_1;
  wire [15:0] Product2_acc_1056_itm_16_1_1;
  wire [15:0] Product2_acc_1086_itm_16_1_1;
  wire [15:0] Product2_acc_1042_itm_16_1_1;
  wire [15:0] Product2_acc_217_itm_17_2_1;
  wire [15:0] Product2_acc_1080_itm_16_1_1;
  wire [15:0] Product2_acc_691_itm_19_4_1;
  wire [15:0] Product2_acc_952_itm_19_4_1;
  wire [15:0] Product2_acc_802_itm_17_2_1;
  wire [15:0] Product2_acc_871_itm_17_2_1;
  wire [15:0] Product2_acc_122_itm_17_2_1;
  wire [15:0] Product2_acc_1144_itm_16_1_1;
  wire [15:0] Product2_acc_733_itm_17_2_1;
  wire [15:0] Product2_acc_216_itm_18_3_1;
  wire [15:0] Product2_acc_285_itm_19_4_1;
  wire [15:0] Product2_acc_531_itm_19_4_1;
  wire [15:0] Product2_acc_299_itm_19_4_1;
  wire [15:0] Product2_acc_450_itm_19_4_1;
  wire [15:0] Product2_acc_1117_itm_16_1_1;
  wire [14:0] Product2_acc_796_itm_18_4_1;
  wire [15:0] Product2_acc_476_itm_19_4_1;
  wire [14:0] Product2_acc_3_itm_15_1_1;
  wire [15:0] Product2_acc_283_itm_18_3_1;
  wire [15:0] Product2_acc_1101_itm_16_1_1;
  wire [15:0] Product2_acc_367_itm_19_4_1;
  wire [15:0] Product2_acc_458_itm_18_3_1;
  wire [15:0] Product2_acc_769_itm_19_4_1;
  wire [15:0] Product2_acc_238_itm_17_2_1;
  wire [15:0] Product2_acc_455_itm_19_4_1;
  wire [14:0] Product2_acc_447_itm_15_1_1;
  wire [15:0] Product2_acc_itm_18_3_1;
  wire [15:0] Product2_acc_152_itm_17_2_1;
  wire [15:0] Product2_acc_554_itm_19_4_1;
  wire [15:0] Product2_acc_1105_itm_16_1_1;
  wire [14:0] Product2_acc_85_itm_15_1_1;
  wire [15:0] Product2_acc_1126_itm_16_1_1;
  wire [15:0] Product2_acc_1118_itm_16_1_1;
  wire [15:0] Product2_acc_954_itm_19_4_1;
  wire [14:0] Product2_acc_629_itm_17_3_1;
  wire [15:0] Product2_acc_1053_itm_16_1_1;
  wire [15:0] Product2_acc_1084_itm_17_2_1;
  wire [15:0] Product2_acc_1114_itm_17_2_1;
  wire [15:0] Product2_acc_666_itm_18_3_1;
  wire [15:0] Product2_acc_1028_itm_17_2_1;
  wire [15:0] Product2_acc_772_itm_18_3_1;
  wire [15:0] Product2_acc_379_itm_18_3_1;
  wire [15:0] Product2_acc_166_itm_18_3_1;
  wire [15:0] Product2_acc_330_itm_19_4_1;
  wire [15:0] Product2_acc_541_itm_19_4_1;
  wire [15:0] Product2_acc_456_itm_19_4_1;
  wire [15:0] Product2_acc_809_itm_19_4_1;
  wire [15:0] Product2_acc_671_itm_18_3_1;
  wire [15:0] Product2_acc_1072_itm_17_2_1;
  wire [15:0] Product2_acc_604_itm_18_3_1;
  wire [15:0] Product2_acc_932_itm_19_4_1;
  wire [15:0] Product2_acc_429_itm_18_3_1;
  wire [15:0] Product2_acc_212_itm_18_3_1;
  wire [15:0] Product2_acc_1066_itm_16_1_1;
  wire [15:0] Product2_acc_937_itm_18_3_1;
  wire [15:0] Product2_acc_8_itm_18_3_1;
  wire [15:0] Product2_acc_528_itm_19_4_1;
  wire [15:0] Product2_acc_727_itm_19_4_1;
  wire [15:0] Product2_acc_876_itm_18_3_1;
  wire [15:0] Product2_acc_72_itm_18_3_1;
  wire [15:0] Product2_acc_141_itm_19_4_1;
  wire [15:0] Product2_acc_499_itm_18_3_1;
  wire [15:0] Product2_acc_281_itm_19_4_1;
  wire [15:0] Product2_acc_1095_itm_16_1_1;
  wire [15:0] Product2_acc_1125_itm_16_1_1;
  wire [15:0] Product2_acc_191_itm_19_4_1;
  wire [15:0] Product2_acc_394_itm_17_2_1;
  wire [15:0] Product2_acc_492_itm_17_2_1;
  wire [15:0] Product2_acc_942_itm_17_2_1;
  wire [15:0] Product2_acc_1079_itm_16_1_1;
  wire [15:0] Product2_acc_154_itm_19_4_1;
  wire [15:0] Product2_acc_547_itm_17_2_1;
  wire [15:0] Product2_acc_901_itm_19_4_1;
  wire [14:0] Product2_acc_62_itm_18_4_1;
  wire [15:0] Product2_acc_601_itm_19_4_1;
  wire [14:0] Product2_acc_801_itm_18_4_1;
  wire [15:0] Product2_acc_742_itm_17_2_1;
  wire [15:0] Product2_acc_298_itm_17_2_1;
  wire [15:0] Product2_acc_560_itm_18_3_1;
  wire [15:0] Product2_acc_670_itm_19_4_1;
  wire [15:0] Product2_acc_795_itm_17_2_1;
  wire [15:0] Product2_acc_664_itm_19_4_1;
  wire [15:0] Product2_acc_951_itm_19_4_1;
  wire [15:0] Product2_acc_11_itm_17_2_1;
  wire [15:0] Product2_acc_193_itm_19_4_1;
  wire [15:0] Product2_acc_398_itm_19_4_1;
  wire [14:0] Product2_acc_603_itm_15_1_1;
  wire [15:0] Product2_acc_73_itm_19_4_1;
  wire [15:0] Product2_acc_606_itm_19_4_1;
  wire [15:0] Product2_acc_374_itm_19_4_1;
  wire [14:0] Product2_acc_1330_itm_17_3_1;
  wire [15:0] Product2_acc_1332_itm_17_2_1;
  wire [14:0] Product2_acc_1334_itm_17_3_1;
  wire [15:0] Product2_acc_1336_itm_18_3_1;
  wire [14:0] Product2_acc_1338_itm_17_3_1;
  wire [8:0] Product2_1_acc_235_itm_11_3_1;
  wire [8:0] Product2_1_acc_386_itm_10_2_1;
  wire [8:0] Product2_1_acc_383_itm_10_2_1;
  wire [8:0] Product2_1_acc_385_itm_10_2_1;
  wire [14:0] Product2_acc_1110_itm_16_2_1;
  wire [14:0] Product2_acc_33_itm_15_1_1;
  wire [14:0] Product2_acc_290_itm_15_1_1;
  wire [14:0] Product2_acc_1147_itm_16_2_1;
  wire [14:0] Product2_acc_887_itm_15_1_1;
  wire [14:0] Product2_acc_91_itm_15_1_1;
  wire [14:0] Product2_acc_448_itm_15_1_1;

  wire[14:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_278_nl;
  wire[16:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_278_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_275_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_275_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_270_nl;
  wire[15:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_270_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_242_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_242_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_300_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_300_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_8_nl;
  wire[10:0] Product2_1_acc_340_nl;
  wire[11:0] nl_Product2_1_acc_340_nl;
  wire[10:0] Product2_1_acc_639_nl;
  wire[11:0] nl_Product2_1_acc_639_nl;
  wire[10:0] Product2_1_acc_640_nl;
  wire[11:0] nl_Product2_1_acc_640_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_299_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_299_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_7_nl;
  wire[10:0] Product2_1_acc_637_nl;
  wire[11:0] nl_Product2_1_acc_637_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_301_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_301_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_9_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_302_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_302_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_10_nl;
  wire[13:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_272_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_272_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_268_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_268_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_222_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_222_nl;
  wire[10:0] Product2_1_acc_300_nl;
  wire[11:0] nl_Product2_1_acc_300_nl;
  wire[10:0] Product2_1_acc_627_nl;
  wire[11:0] nl_Product2_1_acc_627_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_221_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_221_nl;
  wire[10:0] Product2_1_acc_628_nl;
  wire[11:0] nl_Product2_1_acc_628_nl;
  wire[10:0] Product2_1_acc_326_nl;
  wire[11:0] nl_Product2_1_acc_326_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_295_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_295_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_296_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_296_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_264_nl;
  wire[16:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_264_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_187_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_187_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_14_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_186_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_186_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_13_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_185_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_185_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_38_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_184_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_184_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_37_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_183_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_183_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_11_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_182_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_182_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_10_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_181_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_181_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_9_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_180_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_180_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_36_nl;
  wire[11:0] Product2_1_acc_229_nl;
  wire[12:0] nl_Product2_1_acc_229_nl;
  wire[11:0] Product2_1_acc_36_nl;
  wire[12:0] nl_Product2_1_acc_36_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_179_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_179_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_35_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_178_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_178_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_8_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_34_nl;
  wire[13:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_271_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_271_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_263_nl;
  wire[15:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_263_nl;
  wire[8:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_199_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_199_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_nl;
  wire[11:0] Product2_1_acc_174_nl;
  wire[12:0] nl_Product2_1_acc_174_nl;
  wire[8:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_198_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_198_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_50_nl;
  wire[8:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_197_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_197_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_49_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_262_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_262_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_297_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_297_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_5_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_298_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_298_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_6_nl;
  wire[10:0] Product2_1_acc_624_nl;
  wire[11:0] nl_Product2_1_acc_624_nl;
  wire[10:0] Product2_1_acc_625_nl;
  wire[11:0] nl_Product2_1_acc_625_nl;
  wire[10:0] Product2_1_acc_629_nl;
  wire[11:0] nl_Product2_1_acc_629_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_274_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_274_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_267_nl;
  wire[12:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_267_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_249_nl;
  wire[12:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_249_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_227_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_227_nl;
  wire[11:0] Product2_1_acc_252_nl;
  wire[12:0] nl_Product2_1_acc_252_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_226_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_226_nl;
  wire[10:0] Product2_1_acc_622_nl;
  wire[11:0] nl_Product2_1_acc_622_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_247_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_247_nl;
  wire[10:0] Product2_1_acc_374_nl;
  wire[11:0] nl_Product2_1_acc_374_nl;
  wire[10:0] Product2_1_acc_631_nl;
  wire[11:0] nl_Product2_1_acc_631_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_258_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_258_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_225_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_225_nl;
  wire[11:0] Product2_1_acc_34_nl;
  wire[12:0] nl_Product2_1_acc_34_nl;
  wire[10:0] Product2_1_acc_623_nl;
  wire[11:0] nl_Product2_1_acc_623_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_223_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_223_nl;
  wire[10:0] Product2_1_acc_297_nl;
  wire[11:0] nl_Product2_1_acc_297_nl;
  wire[10:0] Product2_1_acc_626_nl;
  wire[11:0] nl_Product2_1_acc_626_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_233_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_233_nl;
  wire[8:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_206_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_206_nl;
  wire[11:0] Product2_1_acc_86_nl;
  wire[12:0] nl_Product2_1_acc_86_nl;
  wire[8:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_205_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_205_nl;
  wire[11:0] Product2_1_acc_104_nl;
  wire[12:0] nl_Product2_1_acc_104_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_228_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_228_nl;
  wire[8:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_196_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_196_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_48_nl;
  wire[10:0] Product2_1_acc_621_nl;
  wire[11:0] nl_Product2_1_acc_621_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_273_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_273_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_265_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_265_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_256_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_256_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_219_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_219_nl;
  wire[10:0] Product2_1_acc_630_nl;
  wire[11:0] nl_Product2_1_acc_630_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_303_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_303_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_254_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_254_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_191_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_191_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_168_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_168_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_51_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_167_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_167_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_52_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_17_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_190_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_190_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_166_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_166_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_53_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_165_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_165_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_21_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_16_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_195_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_195_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_176_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_176_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_6_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_175_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_175_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_5_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_47_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_194_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_194_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_174_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_174_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_173_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_173_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_30_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_45_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_193_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_193_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_172_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_172_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_28_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_171_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_171_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_3_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_44_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_192_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_192_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_170_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_170_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_2_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_169_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_169_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_1_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_18_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_189_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_189_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_164_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_164_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_20_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_163_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_163_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_23_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_15_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_188_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_188_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_162_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_162_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_24_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_39_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_246_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_246_nl;
  wire[10:0] Product2_1_acc_368_nl;
  wire[11:0] nl_Product2_1_acc_368_nl;
  wire[10:0] Product2_1_acc_632_nl;
  wire[11:0] nl_Product2_1_acc_632_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_244_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_244_nl;
  wire[10:0] Product2_1_acc_635_nl;
  wire[11:0] nl_Product2_1_acc_635_nl;
  wire[10:0] Product2_1_acc_303_nl;
  wire[11:0] nl_Product2_1_acc_303_nl;
  wire[15:0] Product2_1_acc_620_nl;
  wire[18:0] nl_Product2_1_acc_620_nl;
  wire[14:0] Product2_1_acc_618_nl;
  wire[16:0] nl_Product2_1_acc_618_nl;
  wire[13:0] Product2_1_acc_614_nl;
  wire[17:0] nl_Product2_1_acc_614_nl;
  wire[11:0] Product2_1_acc_591_nl;
  wire[13:0] nl_Product2_1_acc_591_nl;
  wire[11:0] Product2_1_acc_558_nl;
  wire[12:0] nl_Product2_1_acc_558_nl;
  wire[9:0] Product2_1_acc_517_nl;
  wire[10:0] nl_Product2_1_acc_517_nl;
  wire[11:0] Product2_1_acc_39_nl;
  wire[12:0] nl_Product2_1_acc_39_nl;
  wire[9:0] Product2_1_acc_515_nl;
  wire[10:0] nl_Product2_1_acc_515_nl;
  wire[10:0] Product2_1_acc_307_nl;
  wire[11:0] nl_Product2_1_acc_307_nl;
  wire[11:0] Product2_1_acc_123_nl;
  wire[12:0] nl_Product2_1_acc_123_nl;
  wire[10:0] Product2_1_acc_655_nl;
  wire[11:0] nl_Product2_1_acc_655_nl;
  wire[11:0] Product2_1_acc_488_nl;
  wire[13:0] nl_Product2_1_acc_488_nl;
  wire[10:0] Product2_1_acc_737_nl;
  wire[11:0] nl_Product2_1_acc_737_nl;
  wire[10:0] Product2_1_acc_742_nl;
  wire[11:0] nl_Product2_1_acc_742_nl;
  wire[11:0] Product2_1_acc_489_nl;
  wire[12:0] nl_Product2_1_acc_489_nl;
  wire[10:0] Product2_1_acc_551_nl;
  wire[11:0] nl_Product2_1_acc_551_nl;
  wire[10:0] Product2_1_acc_372_nl;
  wire[11:0] nl_Product2_1_acc_372_nl;
  wire[10:0] Product2_1_acc_446_nl;
  wire[11:0] nl_Product2_1_acc_446_nl;
  wire[10:0] Product2_1_acc_548_nl;
  wire[11:0] nl_Product2_1_acc_548_nl;
  wire[10:0] Product2_1_acc_449_nl;
  wire[11:0] nl_Product2_1_acc_449_nl;
  wire[10:0] Product2_1_acc_279_nl;
  wire[11:0] nl_Product2_1_acc_279_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_279_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_279_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_280_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_280_nl;
  wire[10:0] Product2_1_acc_648_nl;
  wire[11:0] nl_Product2_1_acc_648_nl;
  wire[9:0] Product2_1_acc_717_nl;
  wire[10:0] nl_Product2_1_acc_717_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_281_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_281_nl;
  wire[10:0] Product2_1_acc_736_nl;
  wire[11:0] nl_Product2_1_acc_736_nl;
  wire[10:0] Product2_1_acc_741_nl;
  wire[11:0] nl_Product2_1_acc_741_nl;
  wire[11:0] Product2_1_acc_481_nl;
  wire[12:0] nl_Product2_1_acc_481_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_282_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_282_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_283_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_283_nl;
  wire[10:0] Product2_1_acc_654_nl;
  wire[11:0] nl_Product2_1_acc_654_nl;
  wire[11:0] Product2_1_acc_486_nl;
  wire[13:0] nl_Product2_1_acc_486_nl;
  wire[12:0] Product2_1_acc_605_nl;
  wire[14:0] nl_Product2_1_acc_605_nl;
  wire[11:0] Product2_1_acc_588_nl;
  wire[12:0] nl_Product2_1_acc_588_nl;
  wire[11:0] Product2_1_acc_538_nl;
  wire[12:0] nl_Product2_1_acc_538_nl;
  wire[12:0] Product2_1_acc_115_nl;
  wire[13:0] nl_Product2_1_acc_115_nl;
  wire[10:0] Product2_1_acc_457_nl;
  wire[11:0] nl_Product2_1_acc_457_nl;
  wire[10:0] Product2_1_acc_535_nl;
  wire[11:0] nl_Product2_1_acc_535_nl;
  wire[13:0] Product2_1_acc_137_nl;
  wire[14:0] nl_Product2_1_acc_137_nl;
  wire[11:0] Product2_1_acc_718_nl;
  wire[12:0] nl_Product2_1_acc_718_nl;
  wire[10:0] Product2_1_acc_460_nl;
  wire[11:0] nl_Product2_1_acc_460_nl;
  wire Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_2_nl;
  wire[11:0] Product2_1_acc_543_nl;
  wire[12:0] nl_Product2_1_acc_543_nl;
  wire[12:0] Product2_1_acc_62_nl;
  wire[13:0] nl_Product2_1_acc_62_nl;
  wire[10:0] Product2_1_acc_453_nl;
  wire[11:0] nl_Product2_1_acc_453_nl;
  wire Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_1_nl;
  wire[11:0] Product2_1_acc_540_nl;
  wire[12:0] nl_Product2_1_acc_540_nl;
  wire[11:0] Product2_1_acc_102_nl;
  wire[12:0] nl_Product2_1_acc_102_nl;
  wire[10:0] Product2_1_acc_456_nl;
  wire[11:0] nl_Product2_1_acc_456_nl;
  wire[12:0] Product2_1_acc_587_nl;
  wire[13:0] nl_Product2_1_acc_587_nl;
  wire[10:0] Product2_1_acc_528_nl;
  wire[11:0] nl_Product2_1_acc_528_nl;
  wire[10:0] Product2_1_acc_352_nl;
  wire[11:0] nl_Product2_1_acc_352_nl;
  wire[10:0] Product2_1_acc_465_nl;
  wire[11:0] nl_Product2_1_acc_465_nl;
  wire[10:0] Product2_1_acc_560_nl;
  wire[13:0] nl_Product2_1_acc_560_nl;
  wire[8:0] Product2_1_acc_503_nl;
  wire[10:0] nl_Product2_1_acc_503_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_19_nl;
  wire[8:0] Product2_1_acc_502_nl;
  wire[10:0] nl_Product2_1_acc_502_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_46_nl;
  wire[7:0] Product2_1_acc_496_nl;
  wire[9:0] nl_Product2_1_acc_496_nl;
  wire[6:0] Product2_1_acc_492_nl;
  wire[8:0] nl_Product2_1_acc_492_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_4_nl;
  wire[6:0] Product2_1_acc_491_nl;
  wire[7:0] nl_Product2_1_acc_491_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_12_nl;
  wire[7:0] Product2_1_acc_495_nl;
  wire[9:0] nl_Product2_1_acc_495_nl;
  wire[7:0] Product2_1_acc_494_nl;
  wire[9:0] nl_Product2_1_acc_494_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_7_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_33_nl;
  wire[11:0] Product2_1_acc_584_nl;
  wire[12:0] nl_Product2_1_acc_584_nl;
  wire[10:0] Product2_1_acc_554_nl;
  wire[11:0] nl_Product2_1_acc_554_nl;
  wire[9:0] Product2_1_acc_501_nl;
  wire[12:0] nl_Product2_1_acc_501_nl;
  wire[10:0] Product2_1_acc_442_nl;
  wire[11:0] nl_Product2_1_acc_442_nl;
  wire[10:0] Product2_1_acc_553_nl;
  wire[11:0] nl_Product2_1_acc_553_nl;
  wire[13:0] Product2_1_acc_264_nl;
  wire[14:0] nl_Product2_1_acc_264_nl;
  wire[11:0] Product2_1_acc_719_nl;
  wire[12:0] nl_Product2_1_acc_719_nl;
  wire[13:0] Product2_1_acc_261_nl;
  wire[14:0] nl_Product2_1_acc_261_nl;
  wire[11:0] Product2_1_acc_720_nl;
  wire[12:0] nl_Product2_1_acc_720_nl;
  wire[13:0] Product2_1_acc_602_nl;
  wire[14:0] nl_Product2_1_acc_602_nl;
  wire[12:0] Product2_1_acc_575_nl;
  wire[13:0] nl_Product2_1_acc_575_nl;
  wire[10:0] Product2_1_acc_530_nl;
  wire[11:0] nl_Product2_1_acc_530_nl;
  wire[13:0] Product2_1_acc_175_nl;
  wire[14:0] nl_Product2_1_acc_175_nl;
  wire[11:0] Product2_1_acc_721_nl;
  wire[12:0] nl_Product2_1_acc_721_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_286_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_286_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_2_nl;
  wire[10:0] Product2_1_acc_529_nl;
  wire[11:0] nl_Product2_1_acc_529_nl;
  wire[13:0] Product2_1_acc_192_nl;
  wire[14:0] nl_Product2_1_acc_192_nl;
  wire[10:0] Product2_1_acc_350_nl;
  wire[11:0] nl_Product2_1_acc_350_nl;
  wire[11:0] Product2_1_acc_586_nl;
  wire[14:0] nl_Product2_1_acc_586_nl;
  wire[11:0] Product2_1_acc_172_nl;
  wire[12:0] nl_Product2_1_acc_172_nl;
  wire[11:0] Product2_1_acc_185_nl;
  wire[12:0] nl_Product2_1_acc_185_nl;
  wire[8:0] Product2_1_acc_500_nl;
  wire[10:0] nl_Product2_1_acc_500_nl;
  wire[8:0] Product2_1_acc_499_nl;
  wire[10:0] nl_Product2_1_acc_499_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_43_nl;
  wire[8:0] Product2_1_acc_498_nl;
  wire[10:0] nl_Product2_1_acc_498_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_40_nl;
  wire[8:0] Product2_1_acc_497_nl;
  wire[10:0] nl_Product2_1_acc_497_nl;
  wire[12:0] Product2_1_acc_187_nl;
  wire[13:0] nl_Product2_1_acc_187_nl;
  wire[11:0] Product2_1_acc_200_nl;
  wire[12:0] nl_Product2_1_acc_200_nl;
  wire[12:0] Product2_1_acc_582_nl;
  wire[13:0] nl_Product2_1_acc_582_nl;
  wire[10:0] Product2_1_acc_549_nl;
  wire[11:0] nl_Product2_1_acc_549_nl;
  wire[13:0] Product2_1_acc_7_nl;
  wire[14:0] nl_Product2_1_acc_7_nl;
  wire[10:0] Product2_1_acc_276_nl;
  wire[11:0] nl_Product2_1_acc_276_nl;
  wire[10:0] Product2_1_acc_547_nl;
  wire[11:0] nl_Product2_1_acc_547_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_284_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_284_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_nl;
  wire[10:0] Product2_1_acc_281_nl;
  wire[11:0] nl_Product2_1_acc_281_nl;
  wire[12:0] Product2_1_acc_576_nl;
  wire[13:0] nl_Product2_1_acc_576_nl;
  wire[10:0] Product2_1_acc_532_nl;
  wire[11:0] nl_Product2_1_acc_532_nl;
  wire[11:0] Product2_1_acc_158_nl;
  wire[12:0] nl_Product2_1_acc_158_nl;
  wire[11:0] Product2_1_acc_161_nl;
  wire[12:0] nl_Product2_1_acc_161_nl;
  wire[10:0] Product2_1_acc_531_nl;
  wire[11:0] nl_Product2_1_acc_531_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_285_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_285_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_1_nl;
  wire[10:0] Product2_1_acc_338_nl;
  wire[11:0] nl_Product2_1_acc_338_nl;
  wire[13:0] Product2_1_acc_600_nl;
  wire[14:0] nl_Product2_1_acc_600_nl;
  wire[11:0] Product2_1_acc_581_nl;
  wire[13:0] nl_Product2_1_acc_581_nl;
  wire[11:0] Product2_1_acc_31_nl;
  wire[12:0] nl_Product2_1_acc_31_nl;
  wire[13:0] Product2_1_acc_43_nl;
  wire[14:0] nl_Product2_1_acc_43_nl;
  wire[10:0] Product2_1_acc_289_nl;
  wire[11:0] nl_Product2_1_acc_289_nl;
  wire[11:0] Product2_1_acc_56_nl;
  wire[12:0] nl_Product2_1_acc_56_nl;
  wire[11:0] Product2_1_acc_580_nl;
  wire[12:0] nl_Product2_1_acc_580_nl;
  wire[10:0] Product2_1_acc_544_nl;
  wire[11:0] nl_Product2_1_acc_544_nl;
  wire[11:0] Product2_1_acc_292_nl;
  wire[12:0] nl_Product2_1_acc_292_nl;
  wire[9:0] Product2_1_acc_452_nl;
  wire[10:0] nl_Product2_1_acc_452_nl;
  wire[10:0] Product2_1_acc_293_nl;
  wire[11:0] nl_Product2_1_acc_293_nl;
  wire[10:0] Product2_1_acc_542_nl;
  wire[11:0] nl_Product2_1_acc_542_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_287_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_287_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_3_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_288_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_288_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_4_nl;
  wire[13:0] Product2_1_acc_597_nl;
  wire[14:0] nl_Product2_1_acc_597_nl;
  wire[11:0] Product2_1_acc_573_nl;
  wire[13:0] nl_Product2_1_acc_573_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_nl;
  wire[11:0] Product2_1_acc_572_nl;
  wire[12:0] nl_Product2_1_acc_572_nl;
  wire[10:0] Product2_1_acc_519_nl;
  wire[11:0] nl_Product2_1_acc_519_nl;
  wire[11:0] Product2_1_acc_238_nl;
  wire[12:0] nl_Product2_1_acc_238_nl;
  wire[10:0] Product2_1_acc_518_nl;
  wire[11:0] nl_Product2_1_acc_518_nl;
  wire[10:0] Product2_1_acc_440_nl;
  wire[11:0] nl_Product2_1_acc_440_nl;
  wire[11:0] Product2_1_acc_227_nl;
  wire[12:0] nl_Product2_1_acc_227_nl;
  wire[14:0] Product2_1_acc_619_nl;
  wire[16:0] nl_Product2_1_acc_619_nl;
  wire[14:0] Product2_1_acc_615_nl;
  wire[15:0] nl_Product2_1_acc_615_nl;
  wire[13:0] Product2_1_acc_610_nl;
  wire[18:0] nl_Product2_1_acc_610_nl;
  wire[13:0] Product2_1_acc_258_nl;
  wire[14:0] nl_Product2_1_acc_258_nl;
  wire[13:0] Product2_1_acc_248_nl;
  wire[14:0] nl_Product2_1_acc_248_nl;
  wire[11:0] Product2_1_acc_723_nl;
  wire[12:0] nl_Product2_1_acc_723_nl;
  wire[13:0] Product2_1_acc_231_nl;
  wire[14:0] nl_Product2_1_acc_231_nl;
  wire[11:0] Product2_1_acc_724_nl;
  wire[12:0] nl_Product2_1_acc_724_nl;
  wire[13:0] Product2_1_acc_6_nl;
  wire[14:0] nl_Product2_1_acc_6_nl;
  wire[11:0] Product2_1_acc_725_nl;
  wire[12:0] nl_Product2_1_acc_725_nl;
  wire[11:0] Product2_1_acc_121_nl;
  wire[12:0] nl_Product2_1_acc_121_nl;
  wire[11:0] Product2_1_acc_125_nl;
  wire[12:0] nl_Product2_1_acc_125_nl;
  wire[13:0] Product2_1_acc_126_nl;
  wire[14:0] nl_Product2_1_acc_126_nl;
  wire[11:0] Product2_1_acc_726_nl;
  wire[12:0] nl_Product2_1_acc_726_nl;
  wire[13:0] Product2_1_acc_135_nl;
  wire[14:0] nl_Product2_1_acc_135_nl;
  wire[13:0] Product2_1_acc_94_nl;
  wire[14:0] nl_Product2_1_acc_94_nl;
  wire[11:0] Product2_1_acc_100_nl;
  wire[12:0] nl_Product2_1_acc_100_nl;
  wire[10:0] Product2_1_acc_313_nl;
  wire[11:0] nl_Product2_1_acc_313_nl;
  wire[11:0] Product2_1_acc_111_nl;
  wire[12:0] nl_Product2_1_acc_111_nl;
  wire[13:0] Product2_1_acc_608_nl;
  wire[16:0] nl_Product2_1_acc_608_nl;
  wire[10:0] Product2_1_acc_667_nl;
  wire[11:0] nl_Product2_1_acc_667_nl;
  wire[11:0] Product2_1_acc_472_nl;
  wire[13:0] nl_Product2_1_acc_472_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_292_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_292_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_289_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_289_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_290_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_290_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_291_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_291_nl;
  wire[10:0] Product2_1_acc_666_nl;
  wire[11:0] nl_Product2_1_acc_666_nl;
  wire[9:0] Product2_1_acc_727_nl;
  wire[10:0] nl_Product2_1_acc_727_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_293_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_293_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_294_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_294_nl;
  wire[14:0] Product2_1_acc_609_nl;
  wire[15:0] nl_Product2_1_acc_609_nl;
  wire[12:0] Product2_1_acc_598_nl;
  wire[15:0] nl_Product2_1_acc_598_nl;
  wire[10:0] Product2_1_acc_355_nl;
  wire[11:0] nl_Product2_1_acc_355_nl;
  wire[11:0] Product2_1_acc_213_nl;
  wire[12:0] nl_Product2_1_acc_213_nl;
  wire[11:0] Product2_1_acc_330_nl;
  wire[12:0] nl_Product2_1_acc_330_nl;
  wire[9:0] Product2_1_acc_461_nl;
  wire[10:0] nl_Product2_1_acc_461_nl;
  wire[11:0] Product2_1_acc_151_nl;
  wire[12:0] nl_Product2_1_acc_151_nl;
  wire[10:0] Product2_1_acc_333_nl;
  wire[11:0] nl_Product2_1_acc_333_nl;
  wire[10:0] Product2_1_acc_335_nl;
  wire[11:0] nl_Product2_1_acc_335_nl;
  wire[13:0] Product2_1_acc_215_nl;
  wire[14:0] nl_Product2_1_acc_215_nl;
  wire[12:0] Product2_1_acc_596_nl;
  wire[14:0] nl_Product2_1_acc_596_nl;
  wire[10:0] Product2_1_acc_516_nl;
  wire[11:0] nl_Product2_1_acc_516_nl;
  wire[11:0] Product2_1_acc_46_nl;
  wire[12:0] nl_Product2_1_acc_46_nl;
  wire[9:0] Product2_1_acc_514_nl;
  wire[10:0] nl_Product2_1_acc_514_nl;
  wire[12:0] Product2_1_acc_132_nl;
  wire[13:0] nl_Product2_1_acc_132_nl;
  wire[10:0] Product2_1_acc_513_nl;
  wire[11:0] nl_Product2_1_acc_513_nl;
  wire[11:0] Product2_1_acc_171_nl;
  wire[12:0] nl_Product2_1_acc_171_nl;
  wire[10:0] Product2_1_acc_510_nl;
  wire[11:0] nl_Product2_1_acc_510_nl;
  wire[10:0] Product2_1_acc_441_nl;
  wire[11:0] nl_Product2_1_acc_441_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_27_nl;
  wire[15:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_160_nl;
  wire[16:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_160_nl;
  wire[15:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_157_nl;
  wire[16:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_157_nl;
  wire[14:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_152_nl;
  wire[15:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_152_nl;
  wire[13:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_137_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_137_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_112_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_112_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_111_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_111_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_56_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_56_nl;
  wire[8:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_35_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_35_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_30_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_30_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_32_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_53_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_53_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_144_nl;
  wire[16:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_144_nl;
  wire[12:0] Product2_1_acc_21_nl;
  wire[13:0] nl_Product2_1_acc_21_nl;
  wire[12:0] Product2_1_acc_164_nl;
  wire[13:0] nl_Product2_1_acc_164_nl;
  wire[11:0] Product2_1_acc_168_nl;
  wire[12:0] nl_Product2_1_acc_168_nl;
  wire[12:0] Product2_1_acc_190_nl;
  wire[13:0] nl_Product2_1_acc_190_nl;
  wire[10:0] Product2_1_acc_348_nl;
  wire[11:0] nl_Product2_1_acc_348_nl;
  wire[12:0] Product2_1_acc_218_nl;
  wire[13:0] nl_Product2_1_acc_218_nl;
  wire[13:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_151_nl;
  wire[17:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_151_nl;
  wire[10:0] Product2_1_acc_269_nl;
  wire[11:0] nl_Product2_1_acc_269_nl;
  wire[10:0] Product2_1_acc_274_nl;
  wire[11:0] nl_Product2_1_acc_274_nl;
  wire[12:0] Product2_1_acc_18_nl;
  wire[13:0] nl_Product2_1_acc_18_nl;
  wire[10:0] Product2_1_acc_283_nl;
  wire[11:0] nl_Product2_1_acc_283_nl;
  wire[10:0] Product2_1_acc_286_nl;
  wire[11:0] nl_Product2_1_acc_286_nl;
  wire[10:0] Product2_1_acc_288_nl;
  wire[11:0] nl_Product2_1_acc_288_nl;
  wire[10:0] Product2_1_acc_320_nl;
  wire[11:0] nl_Product2_1_acc_320_nl;
  wire[10:0] Product2_1_acc_322_nl;
  wire[11:0] nl_Product2_1_acc_322_nl;
  wire[10:0] Product2_1_acc_329_nl;
  wire[11:0] nl_Product2_1_acc_329_nl;
  wire[10:0] Product2_1_acc_295_nl;
  wire[11:0] nl_Product2_1_acc_295_nl;
  wire[10:0] Product2_1_acc_302_nl;
  wire[11:0] nl_Product2_1_acc_302_nl;
  wire[10:0] Product2_1_acc_310_nl;
  wire[11:0] nl_Product2_1_acc_310_nl;
  wire[10:0] Product2_1_acc_318_nl;
  wire[11:0] nl_Product2_1_acc_318_nl;
  wire[14:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_156_nl;
  wire[15:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_156_nl;
  wire[13:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_150_nl;
  wire[17:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_150_nl;
  wire[13:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_149_nl;
  wire[16:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_149_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_317_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_317_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_318_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_318_nl;
  wire[10:0] Product2_1_acc_704_nl;
  wire[11:0] nl_Product2_1_acc_704_nl;
  wire[11:0] Product2_1_acc_403_nl;
  wire[13:0] nl_Product2_1_acc_403_nl;
  wire[10:0] Product2_1_acc_705_nl;
  wire[11:0] nl_Product2_1_acc_705_nl;
  wire[11:0] Product2_1_acc_405_nl;
  wire[13:0] nl_Product2_1_acc_405_nl;
  wire[10:0] Product2_1_acc_739_nl;
  wire[11:0] nl_Product2_1_acc_739_nl;
  wire[10:0] Product2_1_acc_744_nl;
  wire[11:0] nl_Product2_1_acc_744_nl;
  wire[11:0] Product2_1_acc_406_nl;
  wire[12:0] nl_Product2_1_acc_406_nl;
  wire[10:0] Product2_1_acc_708_nl;
  wire[11:0] nl_Product2_1_acc_708_nl;
  wire[11:0] Product2_1_acc_409_nl;
  wire[13:0] nl_Product2_1_acc_409_nl;
  wire[10:0] Product2_1_acc_740_nl;
  wire[11:0] nl_Product2_1_acc_740_nl;
  wire[10:0] Product2_1_acc_745_nl;
  wire[11:0] nl_Product2_1_acc_745_nl;
  wire[11:0] Product2_1_acc_412_nl;
  wire[12:0] nl_Product2_1_acc_412_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_319_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_319_nl;
  wire[15:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_159_nl;
  wire[20:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_159_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_22_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_312_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_312_nl;
  wire[10:0] Product2_1_acc_696_nl;
  wire[11:0] nl_Product2_1_acc_696_nl;
  wire[11:0] Product2_1_acc_433_nl;
  wire[13:0] nl_Product2_1_acc_433_nl;
  wire[10:0] Product2_1_acc_687_nl;
  wire[11:0] nl_Product2_1_acc_687_nl;
  wire[11:0] Product2_1_acc_422_nl;
  wire[13:0] nl_Product2_1_acc_422_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_306_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_306_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_307_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_307_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_308_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_308_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_304_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_304_nl;
  wire[10:0] Product2_1_acc_683_nl;
  wire[11:0] nl_Product2_1_acc_683_nl;
  wire[11:0] Product2_1_acc_417_nl;
  wire[13:0] nl_Product2_1_acc_417_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_305_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_305_nl;
  wire[10:0] Product2_1_acc_738_nl;
  wire[11:0] nl_Product2_1_acc_738_nl;
  wire[10:0] Product2_1_acc_743_nl;
  wire[11:0] nl_Product2_1_acc_743_nl;
  wire[10:0] Product2_1_acc_691_nl;
  wire[11:0] nl_Product2_1_acc_691_nl;
  wire[11:0] Product2_1_acc_427_nl;
  wire[13:0] nl_Product2_1_acc_427_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_309_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_309_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_310_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_310_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_311_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_311_nl;
  wire[10:0] Product2_1_acc_697_nl;
  wire[11:0] nl_Product2_1_acc_697_nl;
  wire[11:0] Product2_1_acc_435_nl;
  wire[13:0] nl_Product2_1_acc_435_nl;
  wire[10:0] Product2_1_acc_698_nl;
  wire[11:0] nl_Product2_1_acc_698_nl;
  wire[11:0] Product2_1_acc_437_nl;
  wire[13:0] nl_Product2_1_acc_437_nl;
  wire[13:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_145_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_145_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_119_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_119_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_77_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_77_nl;
  wire[13:0] Product2_1_acc_177_nl;
  wire[14:0] nl_Product2_1_acc_177_nl;
  wire[11:0] Product2_1_acc_729_nl;
  wire[12:0] nl_Product2_1_acc_729_nl;
  wire[11:0] Product2_1_acc_182_nl;
  wire[12:0] nl_Product2_1_acc_182_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_76_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_76_nl;
  wire[10:0] Product2_1_acc_347_nl;
  wire[11:0] nl_Product2_1_acc_347_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_313_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_313_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_11_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_128_nl;
  wire[15:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_128_nl;
  wire[10:0] Product2_1_acc_365_nl;
  wire[11:0] nl_Product2_1_acc_365_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_143_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_143_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_125_nl;
  wire[14:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_125_nl;
  wire[11:0] Product2_1_acc_381_nl;
  wire[12:0] nl_Product2_1_acc_381_nl;
  wire[9:0] Product2_1_acc_387_nl;
  wire[10:0] nl_Product2_1_acc_387_nl;
  wire[13:0] Product2_1_acc_260_nl;
  wire[14:0] nl_Product2_1_acc_260_nl;
  wire[11:0] Product2_1_acc_730_nl;
  wire[12:0] nl_Product2_1_acc_730_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_34_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_34_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_29_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_29_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_31_nl;
  wire[6:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_28_nl;
  wire[8:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_28_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_29_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_124_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_124_nl;
  wire[10:0] Product2_1_acc_390_nl;
  wire[11:0] nl_Product2_1_acc_390_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_314_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_314_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_12_nl;
  wire[10:0] Product2_1_acc_392_nl;
  wire[11:0] nl_Product2_1_acc_392_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_315_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_315_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_13_nl;
  wire[12:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_140_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_140_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_118_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_118_nl;
  wire[10:0] Product2_1_acc_354_nl;
  wire[11:0] nl_Product2_1_acc_354_nl;
  wire[11:0] Product2_1_acc_220_nl;
  wire[12:0] nl_Product2_1_acc_220_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_117_nl;
  wire[13:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_117_nl;
  wire[10:0] Product2_1_acc_397_nl;
  wire[11:0] nl_Product2_1_acc_397_nl;
  wire[10:0] Product2_1_acc_398_nl;
  wire[11:0] nl_Product2_1_acc_398_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_316_nl;
  wire[10:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_316_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_and_14_nl;
  wire[10:0] Product2_1_acc_400_nl;
  wire[11:0] nl_Product2_1_acc_400_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_129_nl;
  wire[12:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_129_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_79_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_79_nl;
  wire[13:0] Product2_1_acc_142_nl;
  wire[14:0] nl_Product2_1_acc_142_nl;
  wire[11:0] Product2_1_acc_728_nl;
  wire[12:0] nl_Product2_1_acc_728_nl;
  wire[11:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_71_nl;
  wire[12:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_71_nl;
  wire[10:0] Product2_1_acc_401_nl;
  wire[11:0] nl_Product2_1_acc_401_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_98_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_98_nl;
  wire[10:0] Product2_1_acc_699_nl;
  wire[11:0] nl_Product2_1_acc_699_nl;
  wire[11:0] Product2_1_acc_439_nl;
  wire[13:0] nl_Product2_1_acc_439_nl;
  wire[9:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_60_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_60_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_33_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_33_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_32_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_32_nl;
  wire[7:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_31_nl;
  wire[9:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_31_nl;
  wire[10:0] nnet_product_mult_layer4_t_config5_weight_t_product_acc_89_nl;
  wire[11:0] nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_89_nl;
  wire[10:0] Product2_1_acc_375_nl;
  wire[11:0] nl_Product2_1_acc_375_nl;
  wire[10:0] Product2_1_acc_389_nl;
  wire[11:0] nl_Product2_1_acc_389_nl;
  wire[15:0] Accum2_acc_220_nl;
  wire[16:0] nl_Accum2_acc_220_nl;
  wire[15:0] Accum2_acc_214_nl;
  wire[17:0] nl_Accum2_acc_214_nl;
  wire[14:0] Accum2_acc_213_nl;
  wire[15:0] nl_Accum2_acc_213_nl;
  wire[7:0] Accum2_acc_1540_nl;
  wire[8:0] nl_Accum2_acc_1540_nl;
  wire[15:0] Accum2_acc_218_nl;
  wire[16:0] nl_Accum2_acc_218_nl;
  wire[15:0] Product2_acc_1233_nl;
  wire[16:0] nl_Product2_acc_1233_nl;
  wire[15:0] Product2_acc_1229_nl;
  wire[16:0] nl_Product2_acc_1229_nl;
  wire[17:0] Product2_acc_1124_nl;
  wire[18:0] nl_Product2_acc_1124_nl;
  wire[15:0] Product2_acc_1222_nl;
  wire[16:0] nl_Product2_acc_1222_nl;
  wire[15:0] Product2_acc_1232_nl;
  wire[17:0] nl_Product2_acc_1232_nl;
  wire[15:0] Product2_acc_1227_nl;
  wire[17:0] nl_Product2_acc_1227_nl;
  wire[14:0] Product2_acc_1224_nl;
  wire[15:0] nl_Product2_acc_1224_nl;
  wire[12:0] Product2_acc_1223_nl;
  wire[13:0] nl_Product2_acc_1223_nl;
  wire[15:0] Accum2_acc_233_nl;
  wire[17:0] nl_Accum2_acc_233_nl;
  wire[15:0] Accum2_acc_230_nl;
  wire[16:0] nl_Accum2_acc_230_nl;
  wire[14:0] Accum2_acc_227_nl;
  wire[16:0] nl_Accum2_acc_227_nl;
  wire[6:0] Accum2_acc_1541_nl;
  wire[7:0] nl_Accum2_acc_1541_nl;
  wire[15:0] Accum2_acc_232_nl;
  wire[17:0] nl_Accum2_acc_232_nl;
  wire[18:0] Product2_acc_530_nl;
  wire[19:0] nl_Product2_acc_530_nl;
  wire[14:0] Product2_acc_1318_nl;
  wire[15:0] Accum2_acc_231_nl;
  wire[16:0] nl_Accum2_acc_231_nl;
  wire[15:0] Accum2_acc_241_nl;
  wire[17:0] nl_Accum2_acc_241_nl;
  wire[5:0] Accum2_acc_1542_nl;
  wire[6:0] nl_Accum2_acc_1542_nl;
  wire[15:0] Accum2_acc_252_nl;
  wire[18:0] nl_Accum2_acc_252_nl;
  wire[4:0] Accum2_acc_1543_nl;
  wire[5:0] nl_Accum2_acc_1543_nl;
  wire[15:0] Accum2_acc_250_nl;
  wire[16:0] nl_Accum2_acc_250_nl;
  wire[15:0] Accum2_acc_249_nl;
  wire[16:0] nl_Accum2_acc_249_nl;
  wire[15:0] Accum2_acc_248_nl;
  wire[16:0] nl_Accum2_acc_248_nl;
  wire[15:0] Accum2_acc_266_nl;
  wire[18:0] nl_Accum2_acc_266_nl;
  wire[15:0] Accum2_acc_265_nl;
  wire[17:0] nl_Accum2_acc_265_nl;
  wire[15:0] Accum2_acc_264_nl;
  wire[17:0] nl_Accum2_acc_264_nl;
  wire[6:0] Accum2_acc_1544_nl;
  wire[7:0] nl_Accum2_acc_1544_nl;
  wire[15:0] Accum2_acc_279_nl;
  wire[17:0] nl_Accum2_acc_279_nl;
  wire[15:0] Accum2_acc_276_nl;
  wire[16:0] nl_Accum2_acc_276_nl;
  wire[14:0] Accum2_acc_272_nl;
  wire[16:0] nl_Accum2_acc_272_nl;
  wire[7:0] Accum2_acc_1545_nl;
  wire[8:0] nl_Accum2_acc_1545_nl;
  wire[15:0] Accum2_acc_278_nl;
  wire[17:0] nl_Accum2_acc_278_nl;
  wire[13:0] Accum2_acc_270_nl;
  wire[14:0] nl_Accum2_acc_270_nl;
  wire[19:0] Product2_acc_369_nl;
  wire[20:0] nl_Product2_acc_369_nl;
  wire[17:0] Product2_acc_1238_nl;
  wire[18:0] nl_Product2_acc_1238_nl;
  wire[12:0] Product2_acc_1319_nl;
  wire[15:0] Accum2_acc_291_nl;
  wire[17:0] nl_Accum2_acc_291_nl;
  wire[15:0] Accum2_acc_287_nl;
  wire[16:0] nl_Accum2_acc_287_nl;
  wire[14:0] Accum2_acc_283_nl;
  wire[15:0] nl_Accum2_acc_283_nl;
  wire[15:0] Accum2_acc_290_nl;
  wire[17:0] nl_Accum2_acc_290_nl;
  wire[15:0] Accum2_acc_289_nl;
  wire[16:0] nl_Accum2_acc_289_nl;
  wire[15:0] Accum2_acc_288_nl;
  wire[16:0] nl_Accum2_acc_288_nl;
  wire[15:0] Accum2_acc_302_nl;
  wire[18:0] nl_Accum2_acc_302_nl;
  wire[6:0] Accum2_acc_1547_nl;
  wire[7:0] nl_Accum2_acc_1547_nl;
  wire[15:0] Accum2_acc_300_nl;
  wire[16:0] nl_Accum2_acc_300_nl;
  wire[15:0] Accum2_acc_314_nl;
  wire[16:0] nl_Accum2_acc_314_nl;
  wire[15:0] Accum2_acc_311_nl;
  wire[17:0] nl_Accum2_acc_311_nl;
  wire[3:0] Accum2_acc_1548_nl;
  wire[4:0] nl_Accum2_acc_1548_nl;
  wire[15:0] Accum2_acc_313_nl;
  wire[16:0] nl_Accum2_acc_313_nl;
  wire[15:0] Accum2_acc_326_nl;
  wire[18:0] nl_Accum2_acc_326_nl;
  wire[12:0] Accum2_acc_317_nl;
  wire[13:0] nl_Accum2_acc_317_nl;
  wire[15:0] Accum2_acc_325_nl;
  wire[16:0] nl_Accum2_acc_325_nl;
  wire[15:0] Accum2_acc_323_nl;
  wire[16:0] nl_Accum2_acc_323_nl;
  wire[14:0] Accum2_acc_320_nl;
  wire[16:0] nl_Accum2_acc_320_nl;
  wire[5:0] Accum2_acc_1549_nl;
  wire[6:0] nl_Accum2_acc_1549_nl;
  wire[15:0] Product2_acc_1248_nl;
  wire[17:0] nl_Product2_acc_1248_nl;
  wire[15:0] Product2_acc_1247_nl;
  wire[18:0] nl_Product2_acc_1247_nl;
  wire[15:0] Product2_acc_1245_nl;
  wire[17:0] nl_Product2_acc_1245_nl;
  wire[15:0] Accum2_acc_338_nl;
  wire[18:0] nl_Accum2_acc_338_nl;
  wire[12:0] Accum2_acc_330_nl;
  wire[13:0] nl_Accum2_acc_330_nl;
  wire[4:0] Accum2_acc_1550_nl;
  wire[5:0] nl_Accum2_acc_1550_nl;
  wire[15:0] Accum2_acc_350_nl;
  wire[17:0] nl_Accum2_acc_350_nl;
  wire[15:0] Accum2_acc_347_nl;
  wire[17:0] nl_Accum2_acc_347_nl;
  wire[15:0] Accum2_acc_349_nl;
  wire[16:0] nl_Accum2_acc_349_nl;
  wire[15:0] Accum2_acc_345_nl;
  wire[16:0] nl_Accum2_acc_345_nl;
  wire[13:0] Accum2_acc_342_nl;
  wire[14:0] nl_Accum2_acc_342_nl;
  wire[5:0] Accum2_acc_1551_nl;
  wire[6:0] nl_Accum2_acc_1551_nl;
  wire[16:0] Product2_acc_1041_nl;
  wire[17:0] nl_Product2_acc_1041_nl;
  wire[15:0] Accum2_acc_348_nl;
  wire[16:0] nl_Accum2_acc_348_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_174_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_174_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_173_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_173_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_168_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_168_nl;
  wire[12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_166_nl;
  wire[13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_166_nl;
  wire[15:0] Accum2_acc_361_nl;
  wire[17:0] nl_Accum2_acc_361_nl;
  wire[15:0] Accum2_acc_360_nl;
  wire[17:0] nl_Accum2_acc_360_nl;
  wire[13:0] Accum2_acc_353_nl;
  wire[14:0] nl_Accum2_acc_353_nl;
  wire[6:0] Accum2_acc_1552_nl;
  wire[7:0] nl_Accum2_acc_1552_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_186_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_186_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_185_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_185_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_179_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_179_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_184_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_184_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_183_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_183_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_182_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_182_nl;
  wire[14:0] nnet_product_mult_input_t_config2_weight_t_product_acc_178_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_178_nl;
  wire[15:0] Accum2_acc_372_nl;
  wire[17:0] nl_Accum2_acc_372_nl;
  wire[15:0] Accum2_acc_371_nl;
  wire[17:0] nl_Accum2_acc_371_nl;
  wire[13:0] Accum2_acc_364_nl;
  wire[14:0] nl_Accum2_acc_364_nl;
  wire[15:0] Accum2_acc_384_nl;
  wire[18:0] nl_Accum2_acc_384_nl;
  wire[3:0] Accum2_acc_1554_nl;
  wire[4:0] nl_Accum2_acc_1554_nl;
  wire[15:0] Accum2_acc_383_nl;
  wire[16:0] nl_Accum2_acc_383_nl;
  wire[15:0] Accum2_acc_382_nl;
  wire[16:0] nl_Accum2_acc_382_nl;
  wire[14:0] Accum2_acc_379_nl;
  wire[16:0] nl_Accum2_acc_379_nl;
  wire[15:0] Accum2_acc_394_nl;
  wire[16:0] nl_Accum2_acc_394_nl;
  wire[15:0] Accum2_acc_390_nl;
  wire[17:0] nl_Accum2_acc_390_nl;
  wire[15:0] Accum2_acc_391_nl;
  wire[16:0] nl_Accum2_acc_391_nl;
  wire[14:0] Accum2_acc_389_nl;
  wire[15:0] nl_Accum2_acc_389_nl;
  wire[15:0] Accum2_acc_405_nl;
  wire[17:0] nl_Accum2_acc_405_nl;
  wire[8:0] Accum2_acc_1555_nl;
  wire[9:0] nl_Accum2_acc_1555_nl;
  wire[15:0] Accum2_acc_404_nl;
  wire[16:0] nl_Accum2_acc_404_nl;
  wire[15:0] Accum2_acc_403_nl;
  wire[16:0] nl_Accum2_acc_403_nl;
  wire[15:0] Accum2_acc_402_nl;
  wire[16:0] nl_Accum2_acc_402_nl;
  wire[14:0] Accum2_acc_398_nl;
  wire[15:0] nl_Accum2_acc_398_nl;
  wire[15:0] Accum2_acc_418_nl;
  wire[16:0] nl_Accum2_acc_418_nl;
  wire[15:0] Accum2_acc_415_nl;
  wire[16:0] nl_Accum2_acc_415_nl;
  wire[15:0] Accum2_acc_414_nl;
  wire[16:0] nl_Accum2_acc_414_nl;
  wire[15:0] Accum2_acc_417_nl;
  wire[18:0] nl_Accum2_acc_417_nl;
  wire[13:0] Accum2_acc_409_nl;
  wire[14:0] nl_Accum2_acc_409_nl;
  wire[5:0] Accum2_acc_1556_nl;
  wire[6:0] nl_Accum2_acc_1556_nl;
  wire[15:0] Accum2_acc_416_nl;
  wire[16:0] nl_Accum2_acc_416_nl;
  wire[15:0] Accum2_acc_428_nl;
  wire[17:0] nl_Accum2_acc_428_nl;
  wire[13:0] Accum2_acc_421_nl;
  wire[14:0] nl_Accum2_acc_421_nl;
  wire[15:0] Accum2_acc_425_nl;
  wire[16:0] nl_Accum2_acc_425_nl;
  wire[14:0] Accum2_acc_422_nl;
  wire[15:0] nl_Accum2_acc_422_nl;
  wire[7:0] Accum2_acc_1557_nl;
  wire[8:0] nl_Accum2_acc_1557_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_201_nl;
  wire[18:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_201_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_198_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_198_nl;
  wire[14:0] nnet_product_mult_input_t_config2_weight_t_product_acc_195_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_195_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_59_nl;
  wire[12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_191_nl;
  wire[13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_191_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_200_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_200_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_199_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_199_nl;
  wire[15:0] Accum2_acc_441_nl;
  wire[18:0] nl_Accum2_acc_441_nl;
  wire[15:0] Accum2_acc_440_nl;
  wire[17:0] nl_Accum2_acc_440_nl;
  wire[15:0] Accum2_acc_439_nl;
  wire[17:0] nl_Accum2_acc_439_nl;
  wire[15:0] Accum2_acc_452_nl;
  wire[17:0] nl_Accum2_acc_452_nl;
  wire[13:0] Accum2_acc_446_nl;
  wire[15:0] nl_Accum2_acc_446_nl;
  wire[5:0] Accum2_acc_1559_nl;
  wire[6:0] nl_Accum2_acc_1559_nl;
  wire[18:0] Product2_acc_617_nl;
  wire[19:0] nl_Product2_acc_617_nl;
  wire[15:0] Accum2_acc_463_nl;
  wire[18:0] nl_Accum2_acc_463_nl;
  wire[4:0] Accum2_acc_1560_nl;
  wire[5:0] nl_Accum2_acc_1560_nl;
  wire[15:0] Accum2_acc_462_nl;
  wire[16:0] nl_Accum2_acc_462_nl;
  wire[15:0] Accum2_acc_458_nl;
  wire[17:0] nl_Accum2_acc_458_nl;
  wire[15:0] Accum2_acc_461_nl;
  wire[16:0] nl_Accum2_acc_461_nl;
  wire[15:0] Accum2_acc_473_nl;
  wire[17:0] nl_Accum2_acc_473_nl;
  wire[15:0] Accum2_acc_471_nl;
  wire[17:0] nl_Accum2_acc_471_nl;
  wire[6:0] Accum2_acc_1561_nl;
  wire[7:0] nl_Accum2_acc_1561_nl;
  wire[15:0] Accum2_acc_484_nl;
  wire[18:0] nl_Accum2_acc_484_nl;
  wire[6:0] Accum2_acc_1562_nl;
  wire[7:0] nl_Accum2_acc_1562_nl;
  wire[15:0] Accum2_acc_483_nl;
  wire[16:0] nl_Accum2_acc_483_nl;
  wire[15:0] Accum2_acc_482_nl;
  wire[16:0] nl_Accum2_acc_482_nl;
  wire[15:0] Accum2_acc_490_nl;
  wire[16:0] nl_Accum2_acc_490_nl;
  wire[12:0] Accum2_acc_487_nl;
  wire[13:0] nl_Accum2_acc_487_nl;
  wire[6:0] Accum2_acc_1563_nl;
  wire[7:0] nl_Accum2_acc_1563_nl;
  wire[15:0] Accum2_acc_501_nl;
  wire[17:0] nl_Accum2_acc_501_nl;
  wire[15:0] Accum2_acc_498_nl;
  wire[16:0] nl_Accum2_acc_498_nl;
  wire[15:0] Accum2_acc_497_nl;
  wire[17:0] nl_Accum2_acc_497_nl;
  wire[13:0] Accum2_acc_493_nl;
  wire[14:0] nl_Accum2_acc_493_nl;
  wire[6:0] Accum2_acc_1564_nl;
  wire[7:0] nl_Accum2_acc_1564_nl;
  wire[15:0] Accum2_acc_516_nl;
  wire[16:0] nl_Accum2_acc_516_nl;
  wire[15:0] Accum2_acc_513_nl;
  wire[16:0] nl_Accum2_acc_513_nl;
  wire[19:0] Product2_acc_678_nl;
  wire[20:0] nl_Product2_acc_678_nl;
  wire[13:0] Product2_acc_1320_nl;
  wire[15:0] Accum2_acc_512_nl;
  wire[17:0] nl_Accum2_acc_512_nl;
  wire[15:0] Accum2_acc_515_nl;
  wire[18:0] nl_Accum2_acc_515_nl;
  wire[4:0] Accum2_acc_1565_nl;
  wire[5:0] nl_Accum2_acc_1565_nl;
  wire[15:0] Accum2_acc_529_nl;
  wire[18:0] nl_Accum2_acc_529_nl;
  wire[15:0] Accum2_acc_528_nl;
  wire[18:0] nl_Accum2_acc_528_nl;
  wire[7:0] Accum2_acc_1566_nl;
  wire[8:0] nl_Accum2_acc_1566_nl;
  wire[13:0] Accum2_acc_536_nl;
  wire[14:0] nl_Accum2_acc_536_nl;
  wire[6:0] Accum2_acc_1567_nl;
  wire[7:0] nl_Accum2_acc_1567_nl;
  wire[15:0] Accum2_acc_552_nl;
  wire[18:0] nl_Accum2_acc_552_nl;
  wire[15:0] Accum2_acc_562_nl;
  wire[16:0] nl_Accum2_acc_562_nl;
  wire[15:0] Accum2_acc_559_nl;
  wire[16:0] nl_Accum2_acc_559_nl;
  wire[19:0] Product2_acc_747_nl;
  wire[20:0] nl_Product2_acc_747_nl;
  wire[17:0] Product2_acc_1253_nl;
  wire[18:0] nl_Product2_acc_1253_nl;
  wire[12:0] Product2_acc_1321_nl;
  wire[15:0] Accum2_acc_558_nl;
  wire[16:0] nl_Accum2_acc_558_nl;
  wire[17:0] Product2_acc_1146_nl;
  wire[18:0] nl_Product2_acc_1146_nl;
  wire[15:0] Product2_acc_1254_nl;
  wire[16:0] nl_Product2_acc_1254_nl;
  wire[15:0] Accum2_acc_561_nl;
  wire[18:0] nl_Accum2_acc_561_nl;
  wire[14:0] Accum2_acc_555_nl;
  wire[16:0] nl_Accum2_acc_555_nl;
  wire[15:0] Accum2_acc_560_nl;
  wire[16:0] nl_Accum2_acc_560_nl;
  wire[15:0] Accum2_acc_574_nl;
  wire[18:0] nl_Accum2_acc_574_nl;
  wire[14:0] Accum2_acc_568_nl;
  wire[16:0] nl_Accum2_acc_568_nl;
  wire[5:0] Accum2_acc_1569_nl;
  wire[6:0] nl_Accum2_acc_1569_nl;
  wire[15:0] Accum2_acc_573_nl;
  wire[17:0] nl_Accum2_acc_573_nl;
  wire[15:0] Accum2_acc_572_nl;
  wire[16:0] nl_Accum2_acc_572_nl;
  wire[16:0] Product2_acc_1104_nl;
  wire[17:0] nl_Product2_acc_1104_nl;
  wire[15:0] Accum2_acc_585_nl;
  wire[17:0] nl_Accum2_acc_585_nl;
  wire[15:0] Accum2_acc_584_nl;
  wire[16:0] nl_Accum2_acc_584_nl;
  wire[3:0] Accum2_acc_1570_nl;
  wire[4:0] nl_Accum2_acc_1570_nl;
  wire[15:0] Accum2_acc_595_nl;
  wire[17:0] nl_Accum2_acc_595_nl;
  wire[15:0] Accum2_acc_594_nl;
  wire[16:0] nl_Accum2_acc_594_nl;
  wire[14:0] Accum2_acc_589_nl;
  wire[15:0] nl_Accum2_acc_589_nl;
  wire[7:0] Accum2_acc_1571_nl;
  wire[8:0] nl_Accum2_acc_1571_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_213_nl;
  wire[18:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_213_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_212_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_212_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_210_nl;
  wire[18:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_210_nl;
  wire[15:0] Accum2_acc_609_nl;
  wire[17:0] nl_Accum2_acc_609_nl;
  wire[13:0] Accum2_acc_603_nl;
  wire[14:0] nl_Accum2_acc_603_nl;
  wire[12:0] Accum2_acc_600_nl;
  wire[13:0] nl_Accum2_acc_600_nl;
  wire[6:0] Accum2_acc_1572_nl;
  wire[7:0] nl_Accum2_acc_1572_nl;
  wire[15:0] Accum2_acc_622_nl;
  wire[16:0] nl_Accum2_acc_622_nl;
  wire[15:0] Accum2_acc_619_nl;
  wire[16:0] nl_Accum2_acc_619_nl;
  wire[19:0] Product2_acc_78_nl;
  wire[20:0] nl_Product2_acc_78_nl;
  wire[17:0] Product2_acc_1256_nl;
  wire[18:0] nl_Product2_acc_1256_nl;
  wire[12:0] Product2_acc_1322_nl;
  wire[15:0] Accum2_acc_618_nl;
  wire[16:0] nl_Accum2_acc_618_nl;
  wire[15:0] Accum2_acc_620_nl;
  wire[17:0] nl_Accum2_acc_620_nl;
  wire[15:0] Accum2_acc_617_nl;
  wire[16:0] nl_Accum2_acc_617_nl;
  wire[17:0] Product2_acc_1111_nl;
  wire[18:0] nl_Product2_acc_1111_nl;
  wire[15:0] Product2_acc_1257_nl;
  wire[16:0] nl_Product2_acc_1257_nl;
  wire[15:0] Accum2_acc_616_nl;
  wire[16:0] nl_Accum2_acc_616_nl;
  wire[14:0] Accum2_acc_613_nl;
  wire[15:0] nl_Accum2_acc_613_nl;
  wire[13:0] Accum2_acc_612_nl;
  wire[14:0] nl_Accum2_acc_612_nl;
  wire[4:0] Accum2_acc_1573_nl;
  wire[5:0] nl_Accum2_acc_1573_nl;
  wire[15:0] Accum2_acc_633_nl;
  wire[18:0] nl_Accum2_acc_633_nl;
  wire[13:0] Accum2_acc_626_nl;
  wire[14:0] nl_Accum2_acc_626_nl;
  wire[6:0] Accum2_acc_1574_nl;
  wire[7:0] nl_Accum2_acc_1574_nl;
  wire[15:0] Accum2_acc_642_nl;
  wire[16:0] nl_Accum2_acc_642_nl;
  wire[13:0] Accum2_acc_637_nl;
  wire[14:0] nl_Accum2_acc_637_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_226_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_226_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_223_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_223_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_222_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_222_nl;
  wire[14:0] nnet_product_mult_input_t_config2_weight_t_product_acc_219_nl;
  wire[15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_219_nl;
  wire[12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_217_nl;
  wire[13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_217_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_225_nl;
  wire[18:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_225_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_224_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_224_nl;
  wire[15:0] Accum2_acc_652_nl;
  wire[18:0] nl_Accum2_acc_652_nl;
  wire[15:0] Accum2_acc_650_nl;
  wire[16:0] nl_Accum2_acc_650_nl;
  wire[15:0] Accum2_acc_649_nl;
  wire[17:0] nl_Accum2_acc_649_nl;
  wire[7:0] Accum2_acc_1576_nl;
  wire[8:0] nl_Accum2_acc_1576_nl;
  wire[15:0] Accum2_acc_665_nl;
  wire[17:0] nl_Accum2_acc_665_nl;
  wire[15:0] Accum2_acc_664_nl;
  wire[18:0] nl_Accum2_acc_664_nl;
  wire[15:0] Accum2_acc_663_nl;
  wire[17:0] nl_Accum2_acc_663_nl;
  wire[15:0] Accum2_acc_676_nl;
  wire[18:0] nl_Accum2_acc_676_nl;
  wire[15:0] Accum2_acc_673_nl;
  wire[16:0] nl_Accum2_acc_673_nl;
  wire[14:0] Accum2_acc_671_nl;
  wire[15:0] nl_Accum2_acc_671_nl;
  wire[13:0] Accum2_acc_669_nl;
  wire[14:0] nl_Accum2_acc_669_nl;
  wire[4:0] Accum2_acc_1578_nl;
  wire[5:0] nl_Accum2_acc_1578_nl;
  wire[15:0] Accum2_acc_674_nl;
  wire[16:0] nl_Accum2_acc_674_nl;
  wire[15:0] Accum2_acc_689_nl;
  wire[16:0] nl_Accum2_acc_689_nl;
  wire[15:0] Accum2_acc_686_nl;
  wire[16:0] nl_Accum2_acc_686_nl;
  wire[15:0] Accum2_acc_685_nl;
  wire[17:0] nl_Accum2_acc_685_nl;
  wire[14:0] Accum2_acc_681_nl;
  wire[15:0] nl_Accum2_acc_681_nl;
  wire[15:0] Accum2_acc_688_nl;
  wire[18:0] nl_Accum2_acc_688_nl;
  wire[5:0] Accum2_acc_1579_nl;
  wire[6:0] nl_Accum2_acc_1579_nl;
  wire[15:0] Accum2_acc_687_nl;
  wire[17:0] nl_Accum2_acc_687_nl;
  wire[15:0] Accum2_acc_700_nl;
  wire[17:0] nl_Accum2_acc_700_nl;
  wire[15:0] Accum2_acc_696_nl;
  wire[17:0] nl_Accum2_acc_696_nl;
  wire[5:0] Accum2_acc_1580_nl;
  wire[6:0] nl_Accum2_acc_1580_nl;
  wire[15:0] Accum2_acc_699_nl;
  wire[17:0] nl_Accum2_acc_699_nl;
  wire[15:0] Accum2_acc_697_nl;
  wire[16:0] nl_Accum2_acc_697_nl;
  wire[19:0] Product2_acc_28_nl;
  wire[20:0] nl_Product2_acc_28_nl;
  wire[13:0] Product2_acc_1323_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_236_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_236_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_235_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_235_nl;
  wire[17:0] Product2_acc_1106_nl;
  wire[18:0] nl_Product2_acc_1106_nl;
  wire[15:0] Product2_acc_1259_nl;
  wire[16:0] nl_Product2_acc_1259_nl;
  wire[13:0] nnet_product_mult_input_t_config2_weight_t_product_acc_230_nl;
  wire[15:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_230_nl;
  wire[15:0] Accum2_acc_713_nl;
  wire[18:0] nl_Accum2_acc_713_nl;
  wire[3:0] Accum2_acc_1581_nl;
  wire[4:0] nl_Accum2_acc_1581_nl;
  wire[15:0] Accum2_acc_712_nl;
  wire[16:0] nl_Accum2_acc_712_nl;
  wire[15:0] Accum2_acc_708_nl;
  wire[16:0] nl_Accum2_acc_708_nl;
  wire[15:0] Accum2_acc_711_nl;
  wire[17:0] nl_Accum2_acc_711_nl;
  wire[15:0] Accum2_acc_724_nl;
  wire[18:0] nl_Accum2_acc_724_nl;
  wire[15:0] Accum2_acc_722_nl;
  wire[16:0] nl_Accum2_acc_722_nl;
  wire[14:0] Accum2_acc_719_nl;
  wire[15:0] nl_Accum2_acc_719_nl;
  wire[4:0] Accum2_acc_1582_nl;
  wire[5:0] nl_Accum2_acc_1582_nl;
  wire[15:0] Accum2_acc_734_nl;
  wire[17:0] nl_Accum2_acc_734_nl;
  wire[15:0] Accum2_acc_733_nl;
  wire[17:0] nl_Accum2_acc_733_nl;
  wire[5:0] Accum2_acc_1583_nl;
  wire[6:0] nl_Accum2_acc_1583_nl;
  wire[15:0] Product2_acc_1270_nl;
  wire[17:0] nl_Product2_acc_1270_nl;
  wire[15:0] Product2_acc_1267_nl;
  wire[17:0] nl_Product2_acc_1267_nl;
  wire[14:0] Product2_acc_1264_nl;
  wire[15:0] nl_Product2_acc_1264_nl;
  wire[15:0] Product2_acc_1269_nl;
  wire[16:0] nl_Product2_acc_1269_nl;
  wire[15:0] Product2_acc_1265_nl;
  wire[17:0] nl_Product2_acc_1265_nl;
  wire[12:0] Product2_acc_1261_nl;
  wire[13:0] nl_Product2_acc_1261_nl;
  wire[12:0] Product2_acc_1260_nl;
  wire[13:0] nl_Product2_acc_1260_nl;
  wire[16:0] Product2_acc_1035_nl;
  wire[17:0] nl_Product2_acc_1035_nl;
  wire[15:0] Accum2_acc_746_nl;
  wire[18:0] nl_Accum2_acc_746_nl;
  wire[15:0] Accum2_acc_745_nl;
  wire[16:0] nl_Accum2_acc_745_nl;
  wire[15:0] Accum2_acc_741_nl;
  wire[16:0] nl_Accum2_acc_741_nl;
  wire[15:0] Accum2_acc_757_nl;
  wire[18:0] nl_Accum2_acc_757_nl;
  wire[12:0] Accum2_acc_749_nl;
  wire[13:0] nl_Accum2_acc_749_nl;
  wire[3:0] Accum2_acc_1585_nl;
  wire[4:0] nl_Accum2_acc_1585_nl;
  wire[15:0] Accum2_acc_755_nl;
  wire[16:0] nl_Accum2_acc_755_nl;
  wire[14:0] Accum2_acc_753_nl;
  wire[16:0] nl_Accum2_acc_753_nl;
  wire[15:0] Accum2_acc_769_nl;
  wire[18:0] nl_Accum2_acc_769_nl;
  wire[19:0] Product2_acc_900_nl;
  wire[20:0] nl_Product2_acc_900_nl;
  wire[15:0] Accum2_acc_768_nl;
  wire[17:0] nl_Accum2_acc_768_nl;
  wire[4:0] Accum2_acc_1586_nl;
  wire[5:0] nl_Accum2_acc_1586_nl;
  wire[15:0] Accum2_acc_779_nl;
  wire[16:0] nl_Accum2_acc_779_nl;
  wire[15:0] Accum2_acc_777_nl;
  wire[18:0] nl_Accum2_acc_777_nl;
  wire[15:0] Accum2_acc_778_nl;
  wire[16:0] nl_Accum2_acc_778_nl;
  wire[15:0] Accum2_acc_787_nl;
  wire[17:0] nl_Accum2_acc_787_nl;
  wire[7:0] Accum2_acc_1588_nl;
  wire[8:0] nl_Accum2_acc_1588_nl;
  wire[15:0] Accum2_acc_786_nl;
  wire[16:0] nl_Accum2_acc_786_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_246_nl;
  wire[18:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_246_nl;
  wire[12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_238_nl;
  wire[13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_238_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_245_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_245_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_244_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_244_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_243_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_243_nl;
  wire[12:0] Accum2_acc_791_nl;
  wire[13:0] nl_Accum2_acc_791_nl;
  wire[6:0] Accum2_acc_1589_nl;
  wire[7:0] nl_Accum2_acc_1589_nl;
  wire[15:0] Accum2_acc_811_nl;
  wire[17:0] nl_Accum2_acc_811_nl;
  wire[4:0] Accum2_acc_1590_nl;
  wire[5:0] nl_Accum2_acc_1590_nl;
  wire[15:0] Accum2_acc_820_nl;
  wire[17:0] nl_Accum2_acc_820_nl;
  wire[15:0] Accum2_acc_818_nl;
  wire[16:0] nl_Accum2_acc_818_nl;
  wire[15:0] Accum2_acc_817_nl;
  wire[16:0] nl_Accum2_acc_817_nl;
  wire[15:0] Accum2_acc_816_nl;
  wire[16:0] nl_Accum2_acc_816_nl;
  wire[15:0] Accum2_acc_833_nl;
  wire[18:0] nl_Accum2_acc_833_nl;
  wire[5:0] Accum2_acc_1591_nl;
  wire[6:0] nl_Accum2_acc_1591_nl;
  wire[15:0] Accum2_acc_844_nl;
  wire[18:0] nl_Accum2_acc_844_nl;
  wire[15:0] Accum2_acc_843_nl;
  wire[16:0] nl_Accum2_acc_843_nl;
  wire[15:0] Accum2_acc_842_nl;
  wire[17:0] nl_Accum2_acc_842_nl;
  wire[13:0] Accum2_acc_837_nl;
  wire[14:0] nl_Accum2_acc_837_nl;
  wire[15:0] Accum2_acc_856_nl;
  wire[18:0] nl_Accum2_acc_856_nl;
  wire[6:0] Accum2_acc_1593_nl;
  wire[7:0] nl_Accum2_acc_1593_nl;
  wire[15:0] Accum2_acc_855_nl;
  wire[17:0] nl_Accum2_acc_855_nl;
  wire[15:0] Accum2_acc_854_nl;
  wire[17:0] nl_Accum2_acc_854_nl;
  wire[15:0] Accum2_acc_867_nl;
  wire[16:0] nl_Accum2_acc_867_nl;
  wire[15:0] Accum2_acc_863_nl;
  wire[17:0] nl_Accum2_acc_863_nl;
  wire[6:0] Accum2_acc_1594_nl;
  wire[7:0] nl_Accum2_acc_1594_nl;
  wire[14:0] Accum2_acc_862_nl;
  wire[16:0] nl_Accum2_acc_862_nl;
  wire[15:0] Accum2_acc_880_nl;
  wire[17:0] nl_Accum2_acc_880_nl;
  wire[15:0] Accum2_acc_876_nl;
  wire[17:0] nl_Accum2_acc_876_nl;
  wire[6:0] Accum2_acc_1595_nl;
  wire[7:0] nl_Accum2_acc_1595_nl;
  wire[15:0] Accum2_acc_879_nl;
  wire[17:0] nl_Accum2_acc_879_nl;
  wire[15:0] Accum2_acc_878_nl;
  wire[16:0] nl_Accum2_acc_878_nl;
  wire[15:0] Accum2_acc_877_nl;
  wire[16:0] nl_Accum2_acc_877_nl;
  wire[15:0] Accum2_acc_893_nl;
  wire[18:0] nl_Accum2_acc_893_nl;
  wire[15:0] Accum2_acc_892_nl;
  wire[16:0] nl_Accum2_acc_892_nl;
  wire[15:0] Accum2_acc_890_nl;
  wire[18:0] nl_Accum2_acc_890_nl;
  wire[6:0] Accum2_acc_1596_nl;
  wire[7:0] nl_Accum2_acc_1596_nl;
  wire[15:0] Accum2_acc_905_nl;
  wire[17:0] nl_Accum2_acc_905_nl;
  wire[15:0] Accum2_acc_904_nl;
  wire[16:0] nl_Accum2_acc_904_nl;
  wire[15:0] Accum2_acc_898_nl;
  wire[16:0] nl_Accum2_acc_898_nl;
  wire[7:0] Accum2_acc_1597_nl;
  wire[8:0] nl_Accum2_acc_1597_nl;
  wire[19:0] Product2_acc_157_nl;
  wire[20:0] nl_Product2_acc_157_nl;
  wire[17:0] Product2_acc_1273_nl;
  wire[18:0] nl_Product2_acc_1273_nl;
  wire[12:0] Product2_acc_1324_nl;
  wire[15:0] Accum2_acc_902_nl;
  wire[16:0] nl_Accum2_acc_902_nl;
  wire[15:0] Accum2_acc_901_nl;
  wire[17:0] nl_Accum2_acc_901_nl;
  wire[15:0] Accum2_acc_916_nl;
  wire[16:0] nl_Accum2_acc_916_nl;
  wire[15:0] Accum2_acc_913_nl;
  wire[16:0] nl_Accum2_acc_913_nl;
  wire[15:0] Accum2_acc_915_nl;
  wire[17:0] nl_Accum2_acc_915_nl;
  wire[13:0] Accum2_acc_910_nl;
  wire[14:0] nl_Accum2_acc_910_nl;
  wire[15:0] Accum2_acc_928_nl;
  wire[18:0] nl_Accum2_acc_928_nl;
  wire[5:0] Accum2_acc_1599_nl;
  wire[6:0] nl_Accum2_acc_1599_nl;
  wire[15:0] Accum2_acc_926_nl;
  wire[16:0] nl_Accum2_acc_926_nl;
  wire[15:0] Accum2_acc_925_nl;
  wire[16:0] nl_Accum2_acc_925_nl;
  wire[15:0] Accum2_acc_940_nl;
  wire[18:0] nl_Accum2_acc_940_nl;
  wire[13:0] Accum2_acc_933_nl;
  wire[14:0] nl_Accum2_acc_933_nl;
  wire[15:0] Accum2_acc_938_nl;
  wire[16:0] nl_Accum2_acc_938_nl;
  wire[14:0] Accum2_acc_935_nl;
  wire[16:0] nl_Accum2_acc_935_nl;
  wire[13:0] Accum2_acc_944_nl;
  wire[14:0] nl_Accum2_acc_944_nl;
  wire[6:0] Accum2_acc_1601_nl;
  wire[7:0] nl_Accum2_acc_1601_nl;
  wire[15:0] Accum2_acc_964_nl;
  wire[17:0] nl_Accum2_acc_964_nl;
  wire[15:0] Accum2_acc_961_nl;
  wire[16:0] nl_Accum2_acc_961_nl;
  wire[14:0] Accum2_acc_958_nl;
  wire[16:0] nl_Accum2_acc_958_nl;
  wire[5:0] Accum2_acc_1602_nl;
  wire[6:0] nl_Accum2_acc_1602_nl;
  wire[15:0] Accum2_acc_963_nl;
  wire[17:0] nl_Accum2_acc_963_nl;
  wire[15:0] Accum2_acc_976_nl;
  wire[17:0] nl_Accum2_acc_976_nl;
  wire[15:0] Accum2_acc_973_nl;
  wire[17:0] nl_Accum2_acc_973_nl;
  wire[15:0] Accum2_acc_975_nl;
  wire[17:0] nl_Accum2_acc_975_nl;
  wire[15:0] Accum2_acc_974_nl;
  wire[17:0] nl_Accum2_acc_974_nl;
  wire[7:0] Accum2_acc_1603_nl;
  wire[8:0] nl_Accum2_acc_1603_nl;
  wire[15:0] Accum2_acc_988_nl;
  wire[17:0] nl_Accum2_acc_988_nl;
  wire[13:0] Accum2_acc_981_nl;
  wire[14:0] nl_Accum2_acc_981_nl;
  wire[12:0] Accum2_acc_979_nl;
  wire[13:0] nl_Accum2_acc_979_nl;
  wire[15:0] Accum2_acc_1000_nl;
  wire[17:0] nl_Accum2_acc_1000_nl;
  wire[14:0] Accum2_acc_995_nl;
  wire[15:0] nl_Accum2_acc_995_nl;
  wire[15:0] Accum2_acc_1013_nl;
  wire[17:0] nl_Accum2_acc_1013_nl;
  wire[15:0] Accum2_acc_1012_nl;
  wire[17:0] nl_Accum2_acc_1012_nl;
  wire[19:0] Product2_acc_644_nl;
  wire[20:0] nl_Product2_acc_644_nl;
  wire[13:0] Product2_acc_1325_nl;
  wire[15:0] Accum2_acc_1023_nl;
  wire[18:0] nl_Accum2_acc_1023_nl;
  wire[7:0] Accum2_acc_1606_nl;
  wire[8:0] nl_Accum2_acc_1606_nl;
  wire[15:0] Accum2_acc_1022_nl;
  wire[16:0] nl_Accum2_acc_1022_nl;
  wire[15:0] Accum2_acc_1035_nl;
  wire[16:0] nl_Accum2_acc_1035_nl;
  wire[15:0] Accum2_acc_1033_nl;
  wire[16:0] nl_Accum2_acc_1033_nl;
  wire[15:0] Accum2_acc_1032_nl;
  wire[18:0] nl_Accum2_acc_1032_nl;
  wire[15:0] Accum2_acc_1034_nl;
  wire[16:0] nl_Accum2_acc_1034_nl;
  wire[15:0] Accum2_acc_1031_nl;
  wire[16:0] nl_Accum2_acc_1031_nl;
  wire[15:0] Accum2_acc_1048_nl;
  wire[16:0] nl_Accum2_acc_1048_nl;
  wire[15:0] Accum2_acc_1046_nl;
  wire[16:0] nl_Accum2_acc_1046_nl;
  wire[15:0] Accum2_acc_1045_nl;
  wire[18:0] nl_Accum2_acc_1045_nl;
  wire[13:0] Accum2_acc_1038_nl;
  wire[14:0] nl_Accum2_acc_1038_nl;
  wire[6:0] Accum2_acc_1608_nl;
  wire[7:0] nl_Accum2_acc_1608_nl;
  wire[15:0] Accum2_acc_1058_nl;
  wire[17:0] nl_Accum2_acc_1058_nl;
  wire[14:0] Accum2_acc_1054_nl;
  wire[16:0] nl_Accum2_acc_1054_nl;
  wire[6:0] Accum2_acc_1609_nl;
  wire[7:0] nl_Accum2_acc_1609_nl;
  wire[15:0] Accum2_acc_1071_nl;
  wire[18:0] nl_Accum2_acc_1071_nl;
  wire[15:0] Accum2_acc_1068_nl;
  wire[16:0] nl_Accum2_acc_1068_nl;
  wire[14:0] Accum2_acc_1064_nl;
  wire[16:0] nl_Accum2_acc_1064_nl;
  wire[5:0] Accum2_acc_1610_nl;
  wire[6:0] nl_Accum2_acc_1610_nl;
  wire[15:0] Accum2_acc_1070_nl;
  wire[17:0] nl_Accum2_acc_1070_nl;
  wire[15:0] Accum2_acc_1084_nl;
  wire[16:0] nl_Accum2_acc_1084_nl;
  wire[15:0] Accum2_acc_1081_nl;
  wire[16:0] nl_Accum2_acc_1081_nl;
  wire[19:0] Product2_acc_41_nl;
  wire[20:0] nl_Product2_acc_41_nl;
  wire[17:0] Product2_acc_1276_nl;
  wire[18:0] nl_Product2_acc_1276_nl;
  wire[12:0] Product2_acc_1326_nl;
  wire[15:0] Accum2_acc_1080_nl;
  wire[16:0] nl_Accum2_acc_1080_nl;
  wire[15:0] Accum2_acc_1082_nl;
  wire[17:0] nl_Accum2_acc_1082_nl;
  wire[15:0] Accum2_acc_1078_nl;
  wire[16:0] nl_Accum2_acc_1078_nl;
  wire[14:0] Accum2_acc_1075_nl;
  wire[16:0] nl_Accum2_acc_1075_nl;
  wire[6:0] Accum2_acc_1611_nl;
  wire[7:0] nl_Accum2_acc_1611_nl;
  wire[15:0] Accum2_acc_1095_nl;
  wire[17:0] nl_Accum2_acc_1095_nl;
  wire[6:0] Accum2_acc_1612_nl;
  wire[7:0] nl_Accum2_acc_1612_nl;
  wire[15:0] Accum2_acc_1094_nl;
  wire[17:0] nl_Accum2_acc_1094_nl;
  wire[15:0] Accum2_acc_1093_nl;
  wire[16:0] nl_Accum2_acc_1093_nl;
  wire[15:0] Accum2_acc_1092_nl;
  wire[17:0] nl_Accum2_acc_1092_nl;
  wire[15:0] Accum2_acc_1107_nl;
  wire[18:0] nl_Accum2_acc_1107_nl;
  wire[6:0] Accum2_acc_1613_nl;
  wire[7:0] nl_Accum2_acc_1613_nl;
  wire[6:0] Accum2_acc_1614_nl;
  wire[7:0] nl_Accum2_acc_1614_nl;
  wire[15:0] Accum2_acc_1138_nl;
  wire[18:0] nl_Accum2_acc_1138_nl;
  wire[15:0] Accum2_acc_1137_nl;
  wire[17:0] nl_Accum2_acc_1137_nl;
  wire[13:0] Accum2_acc_1129_nl;
  wire[14:0] nl_Accum2_acc_1129_nl;
  wire[15:0] Accum2_acc_1136_nl;
  wire[16:0] nl_Accum2_acc_1136_nl;
  wire[15:0] Accum2_acc_1135_nl;
  wire[16:0] nl_Accum2_acc_1135_nl;
  wire[14:0] Accum2_acc_1131_nl;
  wire[15:0] nl_Accum2_acc_1131_nl;
  wire[7:0] Accum2_acc_1615_nl;
  wire[8:0] nl_Accum2_acc_1615_nl;
  wire[15:0] Accum2_acc_1148_nl;
  wire[17:0] nl_Accum2_acc_1148_nl;
  wire[6:0] Accum2_acc_1616_nl;
  wire[7:0] nl_Accum2_acc_1616_nl;
  wire[15:0] Accum2_acc_1155_nl;
  wire[16:0] nl_Accum2_acc_1155_nl;
  wire[14:0] Accum2_acc_1153_nl;
  wire[15:0] nl_Accum2_acc_1153_nl;
  wire[6:0] Accum2_acc_1617_nl;
  wire[7:0] nl_Accum2_acc_1617_nl;
  wire[15:0] Accum2_acc_1167_nl;
  wire[18:0] nl_Accum2_acc_1167_nl;
  wire[12:0] Accum2_acc_1159_nl;
  wire[13:0] nl_Accum2_acc_1159_nl;
  wire[6:0] Accum2_acc_1618_nl;
  wire[7:0] nl_Accum2_acc_1618_nl;
  wire[15:0] Accum2_acc_1166_nl;
  wire[16:0] nl_Accum2_acc_1166_nl;
  wire[15:0] Accum2_acc_1164_nl;
  wire[17:0] nl_Accum2_acc_1164_nl;
  wire[15:0] Accum2_acc_1178_nl;
  wire[17:0] nl_Accum2_acc_1178_nl;
  wire[15:0] Accum2_acc_1173_nl;
  wire[17:0] nl_Accum2_acc_1173_nl;
  wire[6:0] Accum2_acc_1619_nl;
  wire[7:0] nl_Accum2_acc_1619_nl;
  wire[15:0] Accum2_acc_1192_nl;
  wire[17:0] nl_Accum2_acc_1192_nl;
  wire[13:0] Accum2_acc_1184_nl;
  wire[14:0] nl_Accum2_acc_1184_nl;
  wire[6:0] Accum2_acc_1620_nl;
  wire[7:0] nl_Accum2_acc_1620_nl;
  wire[15:0] Accum2_acc_1203_nl;
  wire[17:0] nl_Accum2_acc_1203_nl;
  wire[15:0] Accum2_acc_1199_nl;
  wire[18:0] nl_Accum2_acc_1199_nl;
  wire[15:0] Accum2_acc_1201_nl;
  wire[16:0] nl_Accum2_acc_1201_nl;
  wire[17:0] Product2_acc_1050_nl;
  wire[18:0] nl_Product2_acc_1050_nl;
  wire[15:0] Product2_acc_1277_nl;
  wire[16:0] nl_Product2_acc_1277_nl;
  wire[15:0] Accum2_acc_1215_nl;
  wire[17:0] nl_Accum2_acc_1215_nl;
  wire[15:0] Accum2_acc_1214_nl;
  wire[17:0] nl_Accum2_acc_1214_nl;
  wire[5:0] Accum2_acc_1622_nl;
  wire[6:0] nl_Accum2_acc_1622_nl;
  wire[15:0] Accum2_acc_1228_nl;
  wire[17:0] nl_Accum2_acc_1228_nl;
  wire[15:0] Accum2_acc_1225_nl;
  wire[17:0] nl_Accum2_acc_1225_nl;
  wire[13:0] Accum2_acc_1220_nl;
  wire[14:0] nl_Accum2_acc_1220_nl;
  wire[5:0] Accum2_acc_1623_nl;
  wire[6:0] nl_Accum2_acc_1623_nl;
  wire[15:0] Accum2_acc_1227_nl;
  wire[17:0] nl_Accum2_acc_1227_nl;
  wire[15:0] Accum2_acc_1226_nl;
  wire[16:0] nl_Accum2_acc_1226_nl;
  wire[15:0] Accum2_acc_1240_nl;
  wire[16:0] nl_Accum2_acc_1240_nl;
  wire[15:0] Accum2_acc_1237_nl;
  wire[16:0] nl_Accum2_acc_1237_nl;
  wire[19:0] Product2_acc_174_nl;
  wire[20:0] nl_Product2_acc_174_nl;
  wire[13:0] Product2_acc_1327_nl;
  wire[15:0] Accum2_acc_1236_nl;
  wire[16:0] nl_Accum2_acc_1236_nl;
  wire[15:0] Accum2_acc_1238_nl;
  wire[18:0] nl_Accum2_acc_1238_nl;
  wire[5:0] Accum2_acc_1624_nl;
  wire[6:0] nl_Accum2_acc_1624_nl;
  wire[15:0] Accum2_acc_1254_nl;
  wire[16:0] nl_Accum2_acc_1254_nl;
  wire[15:0] Accum2_acc_1252_nl;
  wire[16:0] nl_Accum2_acc_1252_nl;
  wire[15:0] Accum2_acc_1251_nl;
  wire[16:0] nl_Accum2_acc_1251_nl;
  wire[12:0] Accum2_acc_1243_nl;
  wire[13:0] nl_Accum2_acc_1243_nl;
  wire[5:0] Accum2_acc_1625_nl;
  wire[6:0] nl_Accum2_acc_1625_nl;
  wire[15:0] Accum2_acc_1264_nl;
  wire[17:0] nl_Accum2_acc_1264_nl;
  wire[15:0] Accum2_acc_1262_nl;
  wire[17:0] nl_Accum2_acc_1262_nl;
  wire[13:0] Accum2_acc_1258_nl;
  wire[14:0] nl_Accum2_acc_1258_nl;
  wire[15:0] Accum2_acc_1276_nl;
  wire[17:0] nl_Accum2_acc_1276_nl;
  wire[13:0] Accum2_acc_1270_nl;
  wire[14:0] nl_Accum2_acc_1270_nl;
  wire[15:0] Accum2_acc_1288_nl;
  wire[18:0] nl_Accum2_acc_1288_nl;
  wire[6:0] Accum2_acc_1628_nl;
  wire[7:0] nl_Accum2_acc_1628_nl;
  wire[15:0] Accum2_acc_1297_nl;
  wire[17:0] nl_Accum2_acc_1297_nl;
  wire[15:0] Accum2_acc_1296_nl;
  wire[17:0] nl_Accum2_acc_1296_nl;
  wire[15:0] Accum2_acc_1294_nl;
  wire[16:0] nl_Accum2_acc_1294_nl;
  wire[8:0] Accum2_acc_1629_nl;
  wire[9:0] nl_Accum2_acc_1629_nl;
  wire[15:0] Accum2_acc_1308_nl;
  wire[16:0] nl_Accum2_acc_1308_nl;
  wire[15:0] Accum2_acc_1303_nl;
  wire[16:0] nl_Accum2_acc_1303_nl;
  wire[15:0] Accum2_acc_1305_nl;
  wire[16:0] nl_Accum2_acc_1305_nl;
  wire[15:0] Accum2_acc_1304_nl;
  wire[16:0] nl_Accum2_acc_1304_nl;
  wire[14:0] Accum2_acc_1302_nl;
  wire[16:0] nl_Accum2_acc_1302_nl;
  wire[5:0] Accum2_acc_1630_nl;
  wire[6:0] nl_Accum2_acc_1630_nl;
  wire[15:0] Accum2_acc_1322_nl;
  wire[18:0] nl_Accum2_acc_1322_nl;
  wire[6:0] Accum2_acc_1631_nl;
  wire[7:0] nl_Accum2_acc_1631_nl;
  wire[18:0] Product2_acc_918_nl;
  wire[19:0] nl_Product2_acc_918_nl;
  wire[15:0] Accum2_acc_1334_nl;
  wire[16:0] nl_Accum2_acc_1334_nl;
  wire[15:0] Accum2_acc_1331_nl;
  wire[16:0] nl_Accum2_acc_1331_nl;
  wire[17:0] Product2_acc_717_nl;
  wire[18:0] nl_Product2_acc_717_nl;
  wire[16:0] Product2_acc_1280_nl;
  wire[17:0] nl_Product2_acc_1280_nl;
  wire[12:0] Product2_acc_1328_nl;
  wire[13:0] nl_Product2_acc_1328_nl;
  wire[15:0] Accum2_acc_1330_nl;
  wire[16:0] nl_Accum2_acc_1330_nl;
  wire[14:0] Accum2_acc_1327_nl;
  wire[16:0] nl_Accum2_acc_1327_nl;
  wire[15:0] Accum2_acc_1333_nl;
  wire[18:0] nl_Accum2_acc_1333_nl;
  wire[4:0] Accum2_acc_1632_nl;
  wire[5:0] nl_Accum2_acc_1632_nl;
  wire[15:0] Accum2_acc_1332_nl;
  wire[16:0] nl_Accum2_acc_1332_nl;
  wire[6:0] Accum2_acc_1633_nl;
  wire[7:0] nl_Accum2_acc_1633_nl;
  wire[15:0] Accum2_acc_1354_nl;
  wire[18:0] nl_Accum2_acc_1354_nl;
  wire[15:0] Accum2_acc_1353_nl;
  wire[17:0] nl_Accum2_acc_1353_nl;
  wire[15:0] Accum2_acc_1352_nl;
  wire[16:0] nl_Accum2_acc_1352_nl;
  wire[15:0] Accum2_acc_1351_nl;
  wire[17:0] nl_Accum2_acc_1351_nl;
  wire[15:0] Accum2_acc_1366_nl;
  wire[17:0] nl_Accum2_acc_1366_nl;
  wire[15:0] Accum2_acc_1365_nl;
  wire[16:0] nl_Accum2_acc_1365_nl;
  wire[13:0] Accum2_acc_1359_nl;
  wire[14:0] nl_Accum2_acc_1359_nl;
  wire[15:0] Accum2_acc_1378_nl;
  wire[18:0] nl_Accum2_acc_1378_nl;
  wire[12:0] Accum2_acc_1369_nl;
  wire[13:0] nl_Accum2_acc_1369_nl;
  wire[15:0] Accum2_acc_1377_nl;
  wire[16:0] nl_Accum2_acc_1377_nl;
  wire[14:0] Accum2_acc_1373_nl;
  wire[16:0] nl_Accum2_acc_1373_nl;
  wire[4:0] Accum2_acc_1634_nl;
  wire[5:0] nl_Accum2_acc_1634_nl;
  wire[15:0] Accum2_acc_1376_nl;
  wire[17:0] nl_Accum2_acc_1376_nl;
  wire[15:0] Accum2_acc_1389_nl;
  wire[17:0] nl_Accum2_acc_1389_nl;
  wire[15:0] Accum2_acc_1385_nl;
  wire[16:0] nl_Accum2_acc_1385_nl;
  wire[14:0] Accum2_acc_1382_nl;
  wire[16:0] nl_Accum2_acc_1382_nl;
  wire[6:0] Accum2_acc_1635_nl;
  wire[7:0] nl_Accum2_acc_1635_nl;
  wire[15:0] Accum2_acc_1388_nl;
  wire[17:0] nl_Accum2_acc_1388_nl;
  wire[18:0] Product2_acc_182_nl;
  wire[19:0] nl_Product2_acc_182_nl;
  wire[14:0] Product2_acc_1329_nl;
  wire[15:0] Accum2_acc_1387_nl;
  wire[16:0] nl_Accum2_acc_1387_nl;
  wire[19:0] Product2_acc_922_nl;
  wire[20:0] nl_Product2_acc_922_nl;
  wire[18:0] Product2_acc_1282_nl;
  wire[19:0] nl_Product2_acc_1282_nl;
  wire[15:0] Accum2_acc_1399_nl;
  wire[17:0] nl_Accum2_acc_1399_nl;
  wire[6:0] Accum2_acc_1636_nl;
  wire[7:0] nl_Accum2_acc_1636_nl;
  wire[15:0] Accum2_acc_1412_nl;
  wire[18:0] nl_Accum2_acc_1412_nl;
  wire[15:0] Accum2_acc_1411_nl;
  wire[17:0] nl_Accum2_acc_1411_nl;
  wire[13:0] Accum2_acc_1404_nl;
  wire[14:0] nl_Accum2_acc_1404_nl;
  wire[15:0] Accum2_acc_1410_nl;
  wire[16:0] nl_Accum2_acc_1410_nl;
  wire[15:0] Accum2_acc_nl;
  wire[18:0] nl_Accum2_acc_nl;
  wire[6:0] Accum2_acc_1539_nl;
  wire[7:0] nl_Accum2_acc_1539_nl;
  wire[15:0] Accum2_acc_208_nl;
  wire[16:0] nl_Accum2_acc_208_nl;
  wire[14:0] Accum2_acc_204_nl;
  wire[15:0] nl_Accum2_acc_204_nl;
  wire[15:0] Accum2_acc_1424_nl;
  wire[17:0] nl_Accum2_acc_1424_nl;
  wire[15:0] Accum2_acc_1423_nl;
  wire[17:0] nl_Accum2_acc_1423_nl;
  wire[13:0] Accum2_acc_1415_nl;
  wire[14:0] nl_Accum2_acc_1415_nl;
  wire[6:0] Accum2_acc_1638_nl;
  wire[7:0] nl_Accum2_acc_1638_nl;
  wire[15:0] Accum2_acc_1421_nl;
  wire[16:0] nl_Accum2_acc_1421_nl;
  wire[14:0] Accum2_acc_1416_nl;
  wire[15:0] nl_Accum2_acc_1416_nl;
  wire[15:0] Accum2_acc_1437_nl;
  wire[17:0] nl_Accum2_acc_1437_nl;
  wire[15:0] Accum2_acc_1433_nl;
  wire[16:0] nl_Accum2_acc_1433_nl;
  wire[15:0] Accum2_acc_1436_nl;
  wire[18:0] nl_Accum2_acc_1436_nl;
  wire[5:0] Accum2_acc_1639_nl;
  wire[6:0] nl_Accum2_acc_1639_nl;
  wire[15:0] Accum2_acc_1434_nl;
  wire[16:0] nl_Accum2_acc_1434_nl;
  wire[15:0] Accum2_acc_1448_nl;
  wire[16:0] nl_Accum2_acc_1448_nl;
  wire[14:0] Accum2_acc_1446_nl;
  wire[15:0] nl_Accum2_acc_1446_nl;
  wire[15:0] Accum2_acc_1460_nl;
  wire[18:0] nl_Accum2_acc_1460_nl;
  wire[15:0] Accum2_acc_1459_nl;
  wire[16:0] nl_Accum2_acc_1459_nl;
  wire[15:0] Accum2_acc_1458_nl;
  wire[16:0] nl_Accum2_acc_1458_nl;
  wire[15:0] Accum2_acc_1457_nl;
  wire[17:0] nl_Accum2_acc_1457_nl;
  wire[15:0] Accum2_acc_1474_nl;
  wire[16:0] nl_Accum2_acc_1474_nl;
  wire[15:0] Accum2_acc_1471_nl;
  wire[16:0] nl_Accum2_acc_1471_nl;
  wire[15:0] Accum2_acc_1470_nl;
  wire[16:0] nl_Accum2_acc_1470_nl;
  wire[15:0] Accum2_acc_1473_nl;
  wire[18:0] nl_Accum2_acc_1473_nl;
  wire[4:0] Accum2_acc_1642_nl;
  wire[5:0] nl_Accum2_acc_1642_nl;
  wire[15:0] Accum2_acc_1472_nl;
  wire[16:0] nl_Accum2_acc_1472_nl;
  wire[15:0] Accum2_acc_1467_nl;
  wire[17:0] nl_Accum2_acc_1467_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_260_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_260_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_257_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_257_nl;
  wire[12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_249_nl;
  wire[13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_249_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_259_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_259_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_255_nl;
  wire[17:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_255_nl;
  wire[12:0] nnet_product_mult_input_t_config2_weight_t_product_acc_251_nl;
  wire[13:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_251_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_acc_258_nl;
  wire[16:0] nl_nnet_product_mult_input_t_config2_weight_t_product_acc_258_nl;
  wire[15:0] Accum2_acc_1483_nl;
  wire[16:0] nl_Accum2_acc_1483_nl;
  wire[15:0] Accum2_acc_1481_nl;
  wire[16:0] nl_Accum2_acc_1481_nl;
  wire[14:0] Accum1_2_Accum2_123_Accum2_acc_1_nl;
  wire[15:0] nl_Accum1_2_Accum2_123_Accum2_acc_1_nl;
  wire[5:0] Accum2_acc_1643_nl;
  wire[6:0] nl_Accum2_acc_1643_nl;
  wire[15:0] Accum2_acc_1482_nl;
  wire[16:0] nl_Accum2_acc_1482_nl;
  wire[14:0] Accum2_acc_1480_nl;
  wire[16:0] nl_Accum2_acc_1480_nl;
  wire[13:0] Accum2_acc_1479_nl;
  wire[14:0] nl_Accum2_acc_1479_nl;
  wire[12:0] Accum2_acc_1477_nl;
  wire[13:0] nl_Accum2_acc_1477_nl;
  wire[15:0] Accum2_acc_1492_nl;
  wire[18:0] nl_Accum2_acc_1492_nl;
  wire[6:0] Accum2_acc_1644_nl;
  wire[7:0] nl_Accum2_acc_1644_nl;
  wire[15:0] Accum2_acc_1491_nl;
  wire[16:0] nl_Accum2_acc_1491_nl;
  wire[15:0] Accum2_acc_1504_nl;
  wire[17:0] nl_Accum2_acc_1504_nl;
  wire[15:0] Accum2_acc_1501_nl;
  wire[17:0] nl_Accum2_acc_1501_nl;
  wire[13:0] Accum2_acc_1496_nl;
  wire[14:0] nl_Accum2_acc_1496_nl;
  wire[6:0] Accum2_acc_1645_nl;
  wire[7:0] nl_Accum2_acc_1645_nl;
  wire[15:0] Accum2_acc_1503_nl;
  wire[17:0] nl_Accum2_acc_1503_nl;
  wire[15:0] Accum2_acc_1514_nl;
  wire[16:0] nl_Accum2_acc_1514_nl;
  wire[12:0] Accum2_acc_1507_nl;
  wire[13:0] nl_Accum2_acc_1507_nl;
  wire[15:0] Accum2_acc_1525_nl;
  wire[17:0] nl_Accum2_acc_1525_nl;
  wire[12:0] Accum2_acc_1517_nl;
  wire[13:0] nl_Accum2_acc_1517_nl;
  wire[15:0] Accum2_acc_1524_nl;
  wire[16:0] nl_Accum2_acc_1524_nl;
  wire[15:0] Accum2_acc_1537_nl;
  wire[17:0] nl_Accum2_acc_1537_nl;
  wire[15:0] Accum2_acc_1536_nl;
  wire[18:0] nl_Accum2_acc_1536_nl;
  wire[14:0] Accum1_2_Accum2_128_Accum2_acc_1_nl;
  wire[15:0] nl_Accum1_2_Accum2_128_Accum2_acc_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[13:0] Product2_1_acc_415_nl;
  wire[14:0] nl_Product2_1_acc_415_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_418_nl;
  wire[13:0] nl_Product2_1_acc_418_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_423_nl;
  wire[13:0] nl_Product2_1_acc_423_nl;
  wire[13:0] Product2_1_acc_424_nl;
  wire[14:0] nl_Product2_1_acc_424_nl;
  wire[13:0] Product2_1_acc_425_nl;
  wire[14:0] nl_Product2_1_acc_425_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_428_nl;
  wire[13:0] nl_Product2_1_acc_428_nl;
  wire[12:0] Product2_1_acc_429_nl;
  wire[13:0] nl_Product2_1_acc_429_nl;
  wire[13:0] Product2_1_acc_430_nl;
  wire[14:0] nl_Product2_1_acc_430_nl;
  wire[12:0] Product2_1_acc_431_nl;
  wire[13:0] nl_Product2_1_acc_431_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[11:0] Product2_1_acc_67_nl;
  wire[12:0] nl_Product2_1_acc_67_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[10:0] Product2_1_acc_384_nl;
  wire[11:0] nl_Product2_1_acc_384_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_396_nl;
  wire[13:0] nl_Product2_1_acc_396_nl;
  wire[11:0] Product2_1_acc_76_nl;
  wire[12:0] nl_Product2_1_acc_76_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_391_nl;
  wire[13:0] nl_Product2_1_acc_391_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_393_nl;
  wire[13:0] nl_Product2_1_acc_393_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_399_nl;
  wire[13:0] nl_Product2_1_acc_399_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[10:0] Product2_1_acc_478_nl;
  wire[11:0] nl_Product2_1_acc_478_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[11:0] Product2_1_acc_72_nl;
  wire[12:0] nl_Product2_1_acc_72_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[11:0] Product2_1_acc_241_nl;
  wire[12:0] nl_Product2_1_acc_241_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[10:0] Product2_1_acc_469_nl;
  wire[11:0] nl_Product2_1_acc_469_nl;
  wire[11:0] Product2_1_acc_8_nl;
  wire[12:0] nl_Product2_1_acc_8_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[13:0] Product2_1_acc_410_nl;
  wire[14:0] nl_Product2_1_acc_410_nl;
  wire[13:0] Product2_1_acc_411_nl;
  wire[14:0] nl_Product2_1_acc_411_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_414_nl;
  wire[13:0] nl_Product2_1_acc_414_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[13:0] Product2_1_acc_644_nl;
  wire[14:0] nl_Product2_1_acc_644_nl;
  wire[12:0] Product2_1_acc_645_nl;
  wire[13:0] nl_Product2_1_acc_645_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_633_nl;
  wire[13:0] nl_Product2_1_acc_633_nl;
  wire[12:0] Product2_1_acc_634_nl;
  wire[13:0] nl_Product2_1_acc_634_nl;
  wire[12:0] Product2_1_acc_636_nl;
  wire[13:0] nl_Product2_1_acc_636_nl;
  wire[12:0] Product2_1_acc_638_nl;
  wire[13:0] nl_Product2_1_acc_638_nl;
  wire[12:0] Product2_1_acc_641_nl;
  wire[13:0] nl_Product2_1_acc_641_nl;
  wire[12:0] Product2_1_acc_642_nl;
  wire[13:0] nl_Product2_1_acc_642_nl;
  wire[11:0] Product2_1_acc_79_nl;
  wire[12:0] nl_Product2_1_acc_79_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_41_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire nnet_product_mult_layer4_t_config5_weight_t_product_nor_25_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[13:0] Product2_1_acc_643_nl;
  wire[14:0] nl_Product2_1_acc_643_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[13:0] Product2_1_acc_476_nl;
  wire[14:0] nl_Product2_1_acc_476_nl;
  wire[13:0] Product2_1_acc_477_nl;
  wire[14:0] nl_Product2_1_acc_477_nl;
  wire[13:0] Product2_1_acc_480_nl;
  wire[14:0] nl_Product2_1_acc_480_nl;
  wire[13:0] Product2_1_acc_483_nl;
  wire[14:0] nl_Product2_1_acc_483_nl;
  wire[12:0] Product2_1_acc_484_nl;
  wire[13:0] nl_Product2_1_acc_484_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[12:0] Product2_1_acc_450_nl;
  wire[13:0] nl_Product2_1_acc_450_nl;
  wire[12:0] Product2_1_acc_462_nl;
  wire[13:0] nl_Product2_1_acc_462_nl;
  wire[12:0] Product2_1_acc_464_nl;
  wire[13:0] nl_Product2_1_acc_464_nl;
  wire[12:0] Product2_1_acc_454_nl;
  wire[13:0] nl_Product2_1_acc_454_nl;
  wire[12:0] Product2_1_acc_455_nl;
  wire[13:0] nl_Product2_1_acc_455_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[13:0] Product2_1_acc_466_nl;
  wire[14:0] nl_Product2_1_acc_466_nl;
  wire[12:0] Product2_1_acc_467_nl;
  wire[13:0] nl_Product2_1_acc_467_nl;
  wire[13:0] Product2_1_acc_468_nl;
  wire[14:0] nl_Product2_1_acc_468_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[13:0] Product2_1_acc_473_nl;
  wire[14:0] nl_Product2_1_acc_473_nl;
  wire[13:0] Product2_1_acc_474_nl;
  wire[14:0] nl_Product2_1_acc_474_nl;
  wire[12:0] Product2_1_acc_475_nl;
  wire[13:0] nl_Product2_1_acc_475_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] Product2_acc_1027_nl;
  wire[17:0] nl_Product2_acc_1027_nl;
  wire[17:0] Product2_acc_478_nl;
  wire[18:0] nl_Product2_acc_478_nl;
  wire[17:0] Product2_acc_377_nl;
  wire[18:0] nl_Product2_acc_377_nl;
  wire[18:0] Product2_acc_946_nl;
  wire[19:0] nl_Product2_acc_946_nl;
  wire[16:0] Product2_acc_1064_nl;
  wire[17:0] nl_Product2_acc_1064_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_208_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_219_nl;
  wire[16:0] Product2_acc_1134_nl;
  wire[17:0] nl_Product2_acc_1134_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_53_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_85_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_99_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_60_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_167_nl;
  wire[16:0] Product2_acc_1034_nl;
  wire[17:0] nl_Product2_acc_1034_nl;
  wire[17:0] Product2_acc_297_nl;
  wire[18:0] nl_Product2_acc_297_nl;
  wire[19:0] Product2_acc_75_nl;
  wire[20:0] nl_Product2_acc_75_nl;
  wire[18:0] Product2_acc_728_nl;
  wire[19:0] nl_Product2_acc_728_nl;
  wire[14:0] Product2_acc_1307_nl;
  wire[19:0] Product2_acc_834_nl;
  wire[20:0] nl_Product2_acc_834_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_274_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_66_nl;
  wire[17:0] Product2_acc_934_nl;
  wire[18:0] nl_Product2_acc_934_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_287_nl;
  wire[16:0] Product2_acc_1056_nl;
  wire[17:0] nl_Product2_acc_1056_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_1_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_132_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_301_nl;
  wire[16:0] Product2_acc_1086_nl;
  wire[17:0] nl_Product2_acc_1086_nl;
  wire[16:0] Product2_acc_1042_nl;
  wire[17:0] nl_Product2_acc_1042_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_15_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_336_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_74_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_121_nl;
  wire[17:0] Product2_acc_217_nl;
  wire[18:0] nl_Product2_acc_217_nl;
  wire[16:0] Product2_acc_1080_nl;
  wire[17:0] nl_Product2_acc_1080_nl;
  wire[19:0] Product2_acc_691_nl;
  wire[20:0] nl_Product2_acc_691_nl;
  wire[19:0] Product2_acc_952_nl;
  wire[20:0] nl_Product2_acc_952_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_147_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_258_nl;
  wire[17:0] Product2_acc_802_nl;
  wire[18:0] nl_Product2_acc_802_nl;
  wire[17:0] Product2_acc_871_nl;
  wire[18:0] nl_Product2_acc_871_nl;
  wire[17:0] Product2_acc_122_nl;
  wire[18:0] nl_Product2_acc_122_nl;
  wire[16:0] Product2_acc_1144_nl;
  wire[17:0] nl_Product2_acc_1144_nl;
  wire[17:0] Product2_acc_733_nl;
  wire[18:0] nl_Product2_acc_733_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_203_nl;
  wire[18:0] Product2_acc_216_nl;
  wire[19:0] nl_Product2_acc_216_nl;
  wire[19:0] Product2_acc_285_nl;
  wire[20:0] nl_Product2_acc_285_nl;
  wire[13:0] Product2_acc_1291_nl;
  wire[19:0] Product2_acc_531_nl;
  wire[20:0] nl_Product2_acc_531_nl;
  wire[17:0] Product2_acc_1194_nl;
  wire[18:0] nl_Product2_acc_1194_nl;
  wire[12:0] Product2_acc_1302_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_338_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_244_nl;
  wire[19:0] Product2_acc_299_nl;
  wire[20:0] nl_Product2_acc_299_nl;
  wire[18:0] Product2_acc_1175_nl;
  wire[19:0] nl_Product2_acc_1175_nl;
  wire[19:0] Product2_acc_450_nl;
  wire[20:0] nl_Product2_acc_450_nl;
  wire[17:0] Product2_acc_1186_nl;
  wire[18:0] nl_Product2_acc_1186_nl;
  wire[12:0] Product2_acc_1297_nl;
  wire[16:0] Product2_acc_1117_nl;
  wire[17:0] nl_Product2_acc_1117_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_182_nl;
  wire[18:0] Product2_acc_796_nl;
  wire[19:0] nl_Product2_acc_796_nl;
  wire[14:0] Product2_acc_1310_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_42_nl;
  wire[19:0] Product2_acc_476_nl;
  wire[20:0] nl_Product2_acc_476_nl;
  wire[13:0] Product2_acc_1299_nl;
  wire[15:0] Product2_acc_3_nl;
  wire[16:0] nl_Product2_acc_3_nl;
  wire[18:0] Product2_acc_283_nl;
  wire[19:0] nl_Product2_acc_283_nl;
  wire[14:0] Product2_acc_1290_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_254_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_245_nl;
  wire[16:0] Product2_acc_1101_nl;
  wire[17:0] nl_Product2_acc_1101_nl;
  wire[19:0] Product2_acc_367_nl;
  wire[20:0] nl_Product2_acc_367_nl;
  wire[18:0] Product2_acc_458_nl;
  wire[19:0] nl_Product2_acc_458_nl;
  wire[14:0] Product2_acc_1298_nl;
  wire[19:0] Product2_acc_769_nl;
  wire[20:0] nl_Product2_acc_769_nl;
  wire[18:0] Product2_acc_1208_nl;
  wire[19:0] nl_Product2_acc_1208_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_262_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_229_nl;
  wire[17:0] Product2_acc_238_nl;
  wire[18:0] nl_Product2_acc_238_nl;
  wire[16:0] Product2_acc_1170_nl;
  wire[17:0] nl_Product2_acc_1170_nl;
  wire[12:0] Product2_acc_1289_nl;
  wire[13:0] nl_Product2_acc_1289_nl;
  wire[19:0] Product2_acc_455_nl;
  wire[20:0] nl_Product2_acc_455_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_324_nl;
  wire[15:0] Product2_acc_447_nl;
  wire[16:0] nl_Product2_acc_447_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_162_nl;
  wire[18:0] Product2_acc_nl;
  wire[19:0] nl_Product2_acc_nl;
  wire[14:0] Product2_acc_1283_nl;
  wire[17:0] Product2_acc_152_nl;
  wire[18:0] nl_Product2_acc_152_nl;
  wire[16:0] Product2_acc_1165_nl;
  wire[17:0] nl_Product2_acc_1165_nl;
  wire[12:0] Product2_acc_1286_nl;
  wire[13:0] nl_Product2_acc_1286_nl;
  wire[19:0] Product2_acc_554_nl;
  wire[20:0] nl_Product2_acc_554_nl;
  wire[18:0] Product2_acc_1197_nl;
  wire[19:0] nl_Product2_acc_1197_nl;
  wire[16:0] Product2_acc_1105_nl;
  wire[17:0] nl_Product2_acc_1105_nl;
  wire[15:0] Product2_acc_85_nl;
  wire[16:0] nl_Product2_acc_85_nl;
  wire[16:0] Product2_acc_1126_nl;
  wire[17:0] nl_Product2_acc_1126_nl;
  wire[16:0] Product2_acc_1118_nl;
  wire[17:0] nl_Product2_acc_1118_nl;
  wire[19:0] Product2_acc_954_nl;
  wire[20:0] nl_Product2_acc_954_nl;
  wire[18:0] Product2_acc_1221_nl;
  wire[19:0] nl_Product2_acc_1221_nl;
  wire[17:0] Product2_acc_629_nl;
  wire[18:0] nl_Product2_acc_629_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_nl;
  wire[16:0] Product2_acc_1053_nl;
  wire[17:0] nl_Product2_acc_1053_nl;
  wire[17:0] Product2_acc_1084_nl;
  wire[18:0] nl_Product2_acc_1084_nl;
  wire[15:0] Product2_acc_1184_nl;
  wire[16:0] nl_Product2_acc_1184_nl;
  wire[17:0] Product2_acc_1114_nl;
  wire[18:0] nl_Product2_acc_1114_nl;
  wire[15:0] Product2_acc_1205_nl;
  wire[16:0] nl_Product2_acc_1205_nl;
  wire[18:0] Product2_acc_666_nl;
  wire[19:0] nl_Product2_acc_666_nl;
  wire[14:0] Product2_acc_1305_nl;
  wire[17:0] Product2_acc_1028_nl;
  wire[18:0] nl_Product2_acc_1028_nl;
  wire[15:0] Product2_acc_1161_nl;
  wire[16:0] nl_Product2_acc_1161_nl;
  wire[18:0] Product2_acc_772_nl;
  wire[19:0] nl_Product2_acc_772_nl;
  wire[18:0] Product2_acc_379_nl;
  wire[19:0] nl_Product2_acc_379_nl;
  wire[14:0] Product2_acc_1294_nl;
  wire[18:0] Product2_acc_166_nl;
  wire[19:0] nl_Product2_acc_166_nl;
  wire[19:0] Product2_acc_330_nl;
  wire[20:0] nl_Product2_acc_330_nl;
  wire[17:0] Product2_acc_1178_nl;
  wire[18:0] nl_Product2_acc_1178_nl;
  wire[12:0] Product2_acc_1293_nl;
  wire[19:0] Product2_acc_541_nl;
  wire[20:0] nl_Product2_acc_541_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_311_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_231_nl;
  wire[19:0] Product2_acc_456_nl;
  wire[20:0] nl_Product2_acc_456_nl;
  wire[18:0] Product2_acc_1187_nl;
  wire[19:0] nl_Product2_acc_1187_nl;
  wire[19:0] Product2_acc_809_nl;
  wire[20:0] nl_Product2_acc_809_nl;
  wire[13:0] Product2_acc_1311_nl;
  wire[18:0] Product2_acc_671_nl;
  wire[19:0] nl_Product2_acc_671_nl;
  wire[17:0] Product2_acc_1072_nl;
  wire[18:0] nl_Product2_acc_1072_nl;
  wire[15:0] Product2_acc_1176_nl;
  wire[16:0] nl_Product2_acc_1176_nl;
  wire[18:0] Product2_acc_604_nl;
  wire[19:0] nl_Product2_acc_604_nl;
  wire[14:0] Product2_acc_1304_nl;
  wire[19:0] Product2_acc_932_nl;
  wire[20:0] nl_Product2_acc_932_nl;
  wire[13:0] Product2_acc_1314_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_273_nl;
  wire[18:0] Product2_acc_429_nl;
  wire[19:0] nl_Product2_acc_429_nl;
  wire[18:0] Product2_acc_212_nl;
  wire[19:0] nl_Product2_acc_212_nl;
  wire[14:0] Product2_acc_1288_nl;
  wire[16:0] Product2_acc_1066_nl;
  wire[17:0] nl_Product2_acc_1066_nl;
  wire[18:0] Product2_acc_937_nl;
  wire[19:0] nl_Product2_acc_937_nl;
  wire[14:0] Product2_acc_1315_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_261_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_310_nl;
  wire[18:0] Product2_acc_8_nl;
  wire[19:0] nl_Product2_acc_8_nl;
  wire[19:0] Product2_acc_528_nl;
  wire[20:0] nl_Product2_acc_528_nl;
  wire[13:0] Product2_acc_1301_nl;
  wire[19:0] Product2_acc_727_nl;
  wire[20:0] nl_Product2_acc_727_nl;
  wire[18:0] Product2_acc_876_nl;
  wire[19:0] nl_Product2_acc_876_nl;
  wire[14:0] Product2_acc_1312_nl;
  wire[18:0] Product2_acc_72_nl;
  wire[19:0] nl_Product2_acc_72_nl;
  wire[14:0] Product2_acc_1285_nl;
  wire[19:0] Product2_acc_141_nl;
  wire[20:0] nl_Product2_acc_141_nl;
  wire[18:0] Product2_acc_499_nl;
  wire[19:0] nl_Product2_acc_499_nl;
  wire[19:0] Product2_acc_281_nl;
  wire[20:0] nl_Product2_acc_281_nl;
  wire[16:0] Product2_acc_1095_nl;
  wire[17:0] nl_Product2_acc_1095_nl;
  wire[16:0] Product2_acc_1125_nl;
  wire[17:0] nl_Product2_acc_1125_nl;
  wire[19:0] Product2_acc_191_nl;
  wire[20:0] nl_Product2_acc_191_nl;
  wire[17:0] Product2_acc_394_nl;
  wire[18:0] nl_Product2_acc_394_nl;
  wire[16:0] Product2_acc_1182_nl;
  wire[17:0] nl_Product2_acc_1182_nl;
  wire[12:0] Product2_acc_1295_nl;
  wire[13:0] nl_Product2_acc_1295_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_220_nl;
  wire[17:0] Product2_acc_492_nl;
  wire[18:0] nl_Product2_acc_492_nl;
  wire[16:0] Product2_acc_1191_nl;
  wire[17:0] nl_Product2_acc_1191_nl;
  wire[12:0] Product2_acc_1300_nl;
  wire[13:0] nl_Product2_acc_1300_nl;
  wire[17:0] Product2_acc_942_nl;
  wire[18:0] nl_Product2_acc_942_nl;
  wire[16:0] Product2_acc_1218_nl;
  wire[17:0] nl_Product2_acc_1218_nl;
  wire[12:0] Product2_acc_1316_nl;
  wire[13:0] nl_Product2_acc_1316_nl;
  wire[16:0] Product2_acc_1079_nl;
  wire[17:0] nl_Product2_acc_1079_nl;
  wire[19:0] Product2_acc_154_nl;
  wire[20:0] nl_Product2_acc_154_nl;
  wire[18:0] Product2_acc_1166_nl;
  wire[19:0] nl_Product2_acc_1166_nl;
  wire[17:0] Product2_acc_547_nl;
  wire[18:0] nl_Product2_acc_547_nl;
  wire[16:0] Product2_acc_1196_nl;
  wire[17:0] nl_Product2_acc_1196_nl;
  wire[12:0] Product2_acc_1303_nl;
  wire[13:0] nl_Product2_acc_1303_nl;
  wire[19:0] Product2_acc_901_nl;
  wire[20:0] nl_Product2_acc_901_nl;
  wire[13:0] Product2_acc_1313_nl;
  wire[18:0] Product2_acc_62_nl;
  wire[19:0] nl_Product2_acc_62_nl;
  wire[19:0] Product2_acc_601_nl;
  wire[20:0] nl_Product2_acc_601_nl;
  wire[18:0] Product2_acc_801_nl;
  wire[19:0] nl_Product2_acc_801_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_288_nl;
  wire[17:0] Product2_acc_742_nl;
  wire[18:0] nl_Product2_acc_742_nl;
  wire[16:0] Product2_acc_1207_nl;
  wire[17:0] nl_Product2_acc_1207_nl;
  wire[12:0] Product2_acc_1308_nl;
  wire[13:0] nl_Product2_acc_1308_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_183_nl;
  wire[17:0] Product2_acc_298_nl;
  wire[18:0] nl_Product2_acc_298_nl;
  wire[16:0] Product2_acc_1174_nl;
  wire[17:0] nl_Product2_acc_1174_nl;
  wire[12:0] Product2_acc_1292_nl;
  wire[13:0] nl_Product2_acc_1292_nl;
  wire[18:0] Product2_acc_560_nl;
  wire[19:0] nl_Product2_acc_560_nl;
  wire[19:0] Product2_acc_670_nl;
  wire[20:0] nl_Product2_acc_670_nl;
  wire[17:0] Product2_acc_1203_nl;
  wire[18:0] nl_Product2_acc_1203_nl;
  wire[12:0] Product2_acc_1306_nl;
  wire[17:0] Product2_acc_795_nl;
  wire[18:0] nl_Product2_acc_795_nl;
  wire[16:0] Product2_acc_1210_nl;
  wire[17:0] nl_Product2_acc_1210_nl;
  wire[12:0] Product2_acc_1309_nl;
  wire[13:0] nl_Product2_acc_1309_nl;
  wire[19:0] Product2_acc_664_nl;
  wire[20:0] nl_Product2_acc_664_nl;
  wire[18:0] Product2_acc_1200_nl;
  wire[19:0] nl_Product2_acc_1200_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_300_nl;
  wire[19:0] Product2_acc_951_nl;
  wire[20:0] nl_Product2_acc_951_nl;
  wire[17:0] Product2_acc_1220_nl;
  wire[18:0] nl_Product2_acc_1220_nl;
  wire[12:0] Product2_acc_1317_nl;
  wire[17:0] Product2_acc_11_nl;
  wire[18:0] nl_Product2_acc_11_nl;
  wire[16:0] Product2_acc_1160_nl;
  wire[17:0] nl_Product2_acc_1160_nl;
  wire[12:0] Product2_acc_1284_nl;
  wire[13:0] nl_Product2_acc_1284_nl;
  wire[19:0] Product2_acc_193_nl;
  wire[20:0] nl_Product2_acc_193_nl;
  wire[13:0] Product2_acc_1287_nl;
  wire[19:0] Product2_acc_398_nl;
  wire[20:0] nl_Product2_acc_398_nl;
  wire[13:0] Product2_acc_1296_nl;
  wire[15:0] Product2_acc_603_nl;
  wire[16:0] nl_Product2_acc_603_nl;
  wire nnet_product_mult_input_t_config2_weight_t_product_nor_325_nl;
  wire[19:0] Product2_acc_73_nl;
  wire[20:0] nl_Product2_acc_73_nl;
  wire[18:0] Product2_acc_1163_nl;
  wire[19:0] nl_Product2_acc_1163_nl;
  wire[19:0] Product2_acc_606_nl;
  wire[20:0] nl_Product2_acc_606_nl;
  wire[18:0] Product2_acc_1199_nl;
  wire[19:0] nl_Product2_acc_1199_nl;
  wire[19:0] Product2_acc_374_nl;
  wire[20:0] nl_Product2_acc_374_nl;
  wire[18:0] Product2_acc_1179_nl;
  wire[19:0] nl_Product2_acc_1179_nl;
  wire[17:0] Product2_acc_1330_nl;
  wire[18:0] nl_Product2_acc_1330_nl;
  wire[17:0] Product2_acc_1332_nl;
  wire[18:0] nl_Product2_acc_1332_nl;
  wire[17:0] Product2_acc_1334_nl;
  wire[18:0] nl_Product2_acc_1334_nl;
  wire[18:0] Product2_acc_1336_nl;
  wire[19:0] nl_Product2_acc_1336_nl;
  wire[17:0] Product2_acc_1338_nl;
  wire[18:0] nl_Product2_acc_1338_nl;
  wire[11:0] Product2_1_acc_235_nl;
  wire[12:0] nl_Product2_1_acc_235_nl;
  wire[10:0] Product2_1_acc_386_nl;
  wire[11:0] nl_Product2_1_acc_386_nl;
  wire[10:0] Product2_1_acc_383_nl;
  wire[11:0] nl_Product2_1_acc_383_nl;
  wire[10:0] Product2_1_acc_385_nl;
  wire[11:0] nl_Product2_1_acc_385_nl;
  wire Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_nl;
  wire[16:0] Product2_acc_1110_nl;
  wire[17:0] nl_Product2_acc_1110_nl;
  wire[15:0] Product2_acc_33_nl;
  wire[16:0] nl_Product2_acc_33_nl;
  wire[15:0] Product2_acc_290_nl;
  wire[16:0] nl_Product2_acc_290_nl;
  wire[16:0] Product2_acc_1147_nl;
  wire[17:0] nl_Product2_acc_1147_nl;
  wire[15:0] Product2_acc_887_nl;
  wire[16:0] nl_Product2_acc_887_nl;
  wire[15:0] Product2_acc_91_nl;
  wire[16:0] nl_Product2_acc_91_nl;
  wire[15:0] Product2_acc_448_nl;
  wire[16:0] nl_Product2_acc_448_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [47:0] nl_layer6_out_rsci_idat;
  assign nl_layer6_out_rsci_idat = {layer6_out_rsci_idat_47_32 , layer6_out_rsci_idat_31_16
      , ({{1{layer6_out_rsci_idat_14_0[14]}}, layer6_out_rsci_idat_14_0})};
  converterBlock_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd224)) input_1_rsci (
      .dat(input_1_rsc_dat),
      .idat(input_1_rsci_idat)
    );
  converterBlock_ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd48)) layer6_out_rsci (
      .idat(nl_layer6_out_rsci_idat[47:0]),
      .dat(layer6_out_rsc_dat)
    );
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1540_nl = (nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:6])
      + 8'b00001001;
  assign Accum2_acc_1540_nl = nl_Accum2_acc_1540_nl[7:0];
  assign nl_Accum2_acc_213_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15({Accum2_acc_1540_nl , (nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[5:0])});
  assign Accum2_acc_213_nl = nl_Accum2_acc_213_nl[14:0];
  assign nl_Accum2_acc_214_nl = conv_s2s_15_16(Accum2_acc_213_nl) + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2])
      + conv_s2s_14_16(input_1_rsci_idat[95:82]);
  assign Accum2_acc_214_nl = nl_Accum2_acc_214_nl[15:0];
  assign nl_Accum2_acc_220_nl = Accum2_acc_215_cse_1 + Accum2_acc_214_nl;
  assign Accum2_acc_220_nl = nl_Accum2_acc_220_nl[15:0];
  assign nl_Accum2_acc_218_nl = Product2_acc_191_itm_19_4_1 + Product2_acc_1084_itm_17_2_1;
  assign Accum2_acc_218_nl = nl_Accum2_acc_218_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1 = Accum2_acc_220_nl
      + Accum2_acc_218_nl + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_528_itm_19_4_1 + Product2_acc_601_itm_19_4_1 + Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_727_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[14:10]!=5'b00000);
  assign nl_Product2_acc_1222_nl = (~ (input_1_rsci_idat[191:176])) + conv_s2s_14_16(input_1_rsci_idat[191:178]);
  assign Product2_acc_1222_nl = nl_Product2_acc_1222_nl[15:0];
  assign nl_Product2_acc_1124_nl = conv_s2u_16_18(Product2_acc_1222_nl) + ({(input_1_rsci_idat[191:176])
      , 2'b01});
  assign Product2_acc_1124_nl = nl_Product2_acc_1124_nl[17:0];
  assign nl_Product2_acc_1229_nl = Product2_acc_728_itm_18_3_1 + (readslicef_18_16_2(Product2_acc_1124_nl));
  assign Product2_acc_1229_nl = nl_Product2_acc_1229_nl[15:0];
  assign nl_Product2_acc_1233_nl = Product2_acc_1229_nl + Accum2_acc_215_cse_1;
  assign Product2_acc_1233_nl = nl_Product2_acc_1233_nl[15:0];
  assign nl_Product2_acc_1223_nl = conv_s2s_12_13(input_1_rsci_idat[31:20]) + 13'b0001011000001;
  assign Product2_acc_1223_nl = nl_Product2_acc_1223_nl[12:0];
  assign nl_Product2_acc_1224_nl = conv_s2s_14_15(Product2_acc_122_itm_17_2_1[15:2])
      + conv_s2s_13_15(Product2_acc_1223_nl);
  assign Product2_acc_1224_nl = nl_Product2_acc_1224_nl[14:0];
  assign nl_Product2_acc_1227_nl = (~ (input_1_rsci_idat[31:16])) + conv_s2s_15_16(Product2_acc_1224_nl);
  assign Product2_acc_1227_nl = nl_Product2_acc_1227_nl[15:0];
  assign nl_Product2_acc_1232_nl = Product2_acc_1227_nl + conv_s2s_15_16(input_1_rsci_idat[159:145])
      + conv_s2s_15_16(Product2_acc_1095_itm_16_1_1[15:1]);
  assign Product2_acc_1232_nl = nl_Product2_acc_1232_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1 = Product2_acc_1233_nl
      + Product2_acc_1232_nl + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_281_itm_19_4_1 + Product2_acc_601_itm_19_4_1 + conv_s2s_15_16(Product2_acc_447_itm_15_1_1)
      + conv_s2s_15_16(Product2_acc_itm_18_3_1[15:1]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1541_nl = conv_s2s_6_7(input_1_rsci_idat[79:74]) + 7'b1111111;
  assign Accum2_acc_1541_nl = nl_Accum2_acc_1541_nl[6:0];
  assign nl_Accum2_acc_227_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_15({Accum2_acc_1541_nl , (input_1_rsci_idat[73:68])}) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_227_nl = nl_Accum2_acc_227_nl[14:0];
  assign nl_Accum2_acc_230_nl = Product2_acc_794_cse_sva_1 + conv_s2s_15_16(Accum2_acc_227_nl);
  assign Accum2_acc_230_nl = nl_Accum2_acc_230_nl[15:0];
  assign nl_Accum2_acc_233_nl = Accum2_acc_230_nl + conv_s2s_15_16(Product2_acc_603_itm_15_1_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_233_nl = nl_Accum2_acc_233_nl[15:0];
  assign Product2_acc_1318_nl =  -conv_s2s_14_15(input_1_rsci_idat[127:114]);
  assign nl_Product2_acc_530_nl = conv_s2s_17_19({Product2_acc_1318_nl , (~ (input_1_rsci_idat[113:112]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[127:112])) , 2'b01});
  assign Product2_acc_530_nl = nl_Product2_acc_530_nl[18:0];
  assign nl_Accum2_acc_232_nl = Product2_acc_193_itm_19_4_1 + conv_s2s_15_16(Product2_acc_448_itm_15_1_1)
      + conv_s2s_15_16(readslicef_19_15_4(Product2_acc_530_nl));
  assign Accum2_acc_232_nl = nl_Accum2_acc_232_nl[15:0];
  assign nl_Accum2_acc_231_nl = Product2_acc_367_itm_19_4_1 + Product2_acc_1114_itm_17_2_1;
  assign Accum2_acc_231_nl = nl_Accum2_acc_231_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1 = Accum2_acc_233_nl
      + Accum2_acc_232_nl + Accum2_acc_231_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_241_nl = Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1);
  assign Accum2_acc_241_nl = nl_Accum2_acc_241_nl[15:0];
  assign nl_Accum2_acc_1542_nl = conv_s2s_5_6(input_1_rsci_idat[79:75]) + 6'b111011;
  assign Accum2_acc_1542_nl = nl_Accum2_acc_1542_nl[5:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1 = Accum2_acc_241_nl
      + conv_s2s_15_16(Product2_acc_604_itm_18_3_1[15:1]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_124_cse_sva_1[15:1]) + conv_s2s_13_16({Accum2_acc_1542_nl
      , (input_1_rsci_idat[74:68])}) + conv_s2s_13_16(input_1_rsci_idat[15:3]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1543_nl = conv_s2s_4_5(input_1_rsci_idat[159:156]) + 5'b00001;
  assign Accum2_acc_1543_nl = nl_Accum2_acc_1543_nl[4:0];
  assign nl_Accum2_acc_252_nl = conv_s2s_15_16(input_1_rsci_idat[15:1]) + conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_124_cse_sva_1[15:2]) + conv_s2s_13_16({Accum2_acc_1543_nl
      , (input_1_rsci_idat[155:148])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_252_nl = nl_Accum2_acc_252_nl[15:0];
  assign nl_Accum2_acc_250_nl = Product2_acc_368_cse_sva_1 + Product2_acc_450_itm_19_4_1;
  assign Accum2_acc_250_nl = nl_Accum2_acc_250_nl[15:0];
  assign nl_Accum2_acc_249_nl = Product2_acc_531_itm_19_4_1 + Product2_acc_730_cse_sva_1;
  assign Accum2_acc_249_nl = nl_Accum2_acc_249_nl[15:0];
  assign nl_Accum2_acc_248_nl = Product2_acc_795_itm_17_2_1 + Product2_acc_932_itm_19_4_1;
  assign Accum2_acc_248_nl = nl_Accum2_acc_248_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1 = Accum2_acc_252_nl
      + Accum2_acc_250_nl + Product2_acc_191_itm_19_4_1 + Product2_acc_1336_itm_18_3_1
      + Accum2_acc_249_nl + Accum2_acc_248_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_266_nl = conv_s2s_15_16(Product2_acc_796_itm_18_4_1) + conv_s2s_15_16(Product2_acc_867_cse_sva_1[15:1])
      + conv_s2s_14_16(input_1_rsci_idat[143:130]) + conv_s2s_14_16(Product2_acc_447_itm_15_1_1[14:1])
      + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1);
  assign Accum2_acc_266_nl = nl_Accum2_acc_266_nl[15:0];
  assign nl_Accum2_acc_265_nl = Accum2_acc_261_cse_1 + conv_s2s_15_16(Product2_acc_283_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_3_itm_15_1_1);
  assign Accum2_acc_265_nl = nl_Accum2_acc_265_nl[15:0];
  assign nl_Accum2_acc_1544_nl = conv_s2s_6_7(input_1_rsci_idat[47:42]) + 7'b1111111;
  assign Accum2_acc_1544_nl = nl_Accum2_acc_1544_nl[6:0];
  assign nl_Accum2_acc_264_nl = Product2_acc_664_itm_19_4_1 + conv_s2s_15_16(Product2_acc_62_itm_18_4_1)
      + conv_s2s_14_16({Accum2_acc_1544_nl , (input_1_rsci_idat[41:35])});
  assign Accum2_acc_264_nl = nl_Accum2_acc_264_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1 = Accum2_acc_266_nl
      + Accum2_acc_265_nl + Accum2_acc_264_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1545_nl = conv_s2s_7_8(input_1_rsci_idat[111:105]) + 8'b00000001;
  assign Accum2_acc_1545_nl = nl_Accum2_acc_1545_nl[7:0];
  assign nl_Accum2_acc_272_nl = conv_s2s_14_15({Accum2_acc_1545_nl , (input_1_rsci_idat[104:99])})
      + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_15(input_1_rsci_idat[47:35]);
  assign Accum2_acc_272_nl = nl_Accum2_acc_272_nl[14:0];
  assign nl_Accum2_acc_276_nl = Product2_acc_797_cse_sva_1 + conv_s2s_15_16(Accum2_acc_272_nl);
  assign Accum2_acc_276_nl = nl_Accum2_acc_276_nl[15:0];
  assign nl_Accum2_acc_279_nl = Accum2_acc_276_nl + conv_s2s_15_16(input_1_rsci_idat[127:113])
      + conv_s2s_14_16(Product2_acc_934_itm_17_2_1[15:2]) + conv_s2s_14_16(input_1_rsci_idat[143:130]);
  assign Accum2_acc_279_nl = nl_Accum2_acc_279_nl[15:0];
  assign nl_Accum2_acc_270_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign Accum2_acc_270_nl = nl_Accum2_acc_270_nl[13:0];
  assign nl_Accum2_acc_278_nl = conv_s2s_15_16(Product2_acc_733_itm_17_2_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_1332_itm_17_2_1[15:1]) + conv_s2s_14_16(Accum2_acc_270_nl);
  assign Accum2_acc_278_nl = nl_Accum2_acc_278_nl[15:0];
  assign Product2_acc_1319_nl =  -conv_s2s_12_13(input_1_rsci_idat[95:84]);
  assign nl_Product2_acc_1238_nl = ({(input_1_rsci_idat[95:80]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1319_nl
      , (~ (input_1_rsci_idat[83:80]))});
  assign Product2_acc_1238_nl = nl_Product2_acc_1238_nl[17:0];
  assign nl_Product2_acc_369_nl = conv_s2s_18_20(Product2_acc_1238_nl) + ({(~ (input_1_rsci_idat[95:80]))
      , 4'b0000});
  assign Product2_acc_369_nl = nl_Product2_acc_369_nl[19:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1 = Accum2_acc_279_nl
      + Accum2_acc_278_nl + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + (readslicef_20_16_4(Product2_acc_369_nl));
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_283_nl = conv_s2s_14_15(Product2_acc_871_itm_17_2_1[15:2])
      + conv_s2s_13_15({Accum2_Accum2_conc_127_12_7 , (input_1_rsci_idat[170:164])});
  assign Accum2_acc_283_nl = nl_Accum2_acc_283_nl[14:0];
  assign nl_Accum2_acc_287_nl = Product2_acc_1125_itm_16_1_1 + conv_s2s_15_16(Accum2_acc_283_nl);
  assign Accum2_acc_287_nl = nl_Accum2_acc_287_nl[15:0];
  assign nl_Accum2_acc_291_nl = Accum2_acc_287_nl + conv_s2s_15_16(input_1_rsci_idat[223:209])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_291_nl = nl_Accum2_acc_291_nl[15:0];
  assign nl_Accum2_acc_290_nl = Accum2_acc_285_cse_1 + conv_s2s_15_16(Product2_acc_1332_itm_17_2_1[15:1])
      + conv_s2s_13_16(input_1_rsci_idat[127:115]) + conv_s2s_12_16(input_1_rsci_idat[47:36]);
  assign Accum2_acc_290_nl = nl_Accum2_acc_290_nl[15:0];
  assign nl_Accum2_acc_289_nl = Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_1084_itm_17_2_1;
  assign Accum2_acc_289_nl = nl_Accum2_acc_289_nl[15:0];
  assign nl_Accum2_acc_288_nl = Product2_acc_606_itm_19_4_1 + Product2_acc_665_cse_sva_1;
  assign Accum2_acc_288_nl = nl_Accum2_acc_288_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1 = Accum2_acc_291_nl
      + Accum2_acc_290_nl + Accum2_acc_289_nl + Accum2_acc_288_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1547_nl = conv_s2s_6_7(input_1_rsci_idat[47:42]) + 7'b1111101;
  assign Accum2_acc_1547_nl = nl_Accum2_acc_1547_nl[6:0];
  assign nl_Accum2_acc_302_nl = conv_s2s_15_16(Product2_acc_604_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1]) + conv_s2s_14_16(Accum2_acc_295_cse_1)
      + conv_s2s_14_16({Accum2_acc_1547_nl , (input_1_rsci_idat[41:35])}) + conv_s2s_14_16(Product2_acc_733_itm_17_2_1[15:2]);
  assign Accum2_acc_302_nl = nl_Accum2_acc_302_nl[15:0];
  assign nl_Accum2_acc_300_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_532_cse_sva_1;
  assign Accum2_acc_300_nl = nl_Accum2_acc_300_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1 = Accum2_acc_302_nl
      + Accum2_acc_300_nl + Product2_acc_666_itm_18_3_1 + Product2_acc_932_itm_19_4_1
      + Product2_acc_191_itm_19_4_1 + Product2_acc_285_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1548_nl = conv_s2s_3_4(input_1_rsci_idat[191:189]) + 4'b1111;
  assign Accum2_acc_1548_nl = nl_Accum2_acc_1548_nl[3:0];
  assign nl_Accum2_acc_311_nl = conv_s2s_15_16(Product2_acc_447_itm_15_1_1) + conv_s2s_13_16(Accum2_acc_306_cse_1)
      + conv_s2s_13_16({Accum2_acc_1548_nl , (input_1_rsci_idat[188:180])});
  assign Accum2_acc_311_nl = nl_Accum2_acc_311_nl[15:0];
  assign nl_Accum2_acc_314_nl = Accum2_acc_311_nl + Product2_acc_1064_itm_16_1_1;
  assign Accum2_acc_314_nl = nl_Accum2_acc_314_nl[15:0];
  assign nl_Accum2_acc_313_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_936_cse_sva_1;
  assign Accum2_acc_313_nl = nl_Accum2_acc_313_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1 = Accum2_acc_314_nl
      + Accum2_acc_313_nl + conv_s2s_14_16(Product2_acc_532_cse_sva_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[95:83]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_317_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[15:4]);
  assign Accum2_acc_317_nl = nl_Accum2_acc_317_nl[12:0];
  assign nl_Accum2_acc_326_nl = conv_s2s_15_16(Product2_acc_937_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_124_cse_sva_1[15:2]) + conv_s2s_13_16(Accum2_acc_317_nl);
  assign Accum2_acc_326_nl = nl_Accum2_acc_326_nl[15:0];
  assign nl_Accum2_acc_325_nl = Product2_acc_195_cse_sva_1 + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_325_nl = nl_Accum2_acc_325_nl[15:0];
  assign nl_Accum2_acc_1549_nl = conv_s2s_5_6(input_1_rsci_idat[159:155]) + 6'b000011;
  assign Accum2_acc_1549_nl = nl_Accum2_acc_1549_nl[5:0];
  assign nl_Accum2_acc_320_nl = conv_s2s_14_15(input_1_rsci_idat[191:178]) + conv_s2s_13_15({Accum2_acc_1549_nl
      , (input_1_rsci_idat[154:148])}) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign Accum2_acc_320_nl = nl_Accum2_acc_320_nl[14:0];
  assign nl_Accum2_acc_323_nl = Product2_acc_1114_itm_17_2_1 + conv_s2s_15_16(Accum2_acc_320_nl);
  assign Accum2_acc_323_nl = nl_Accum2_acc_323_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1 = Accum2_acc_326_nl
      + Accum2_acc_325_nl + Accum2_acc_323_nl + Product2_acc_455_itm_19_4_1 + Product2_acc_560_itm_18_3_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[14:10]!=5'b00000);
  assign nl_Product2_acc_1248_nl = Accum2_acc_261_cse_1 + conv_s2s_15_16(input_1_rsci_idat[159:145])
      + conv_s2s_15_16(input_1_rsci_idat[191:177]);
  assign Product2_acc_1248_nl = nl_Product2_acc_1248_nl[15:0];
  assign nl_Product2_acc_1247_nl = conv_s2s_15_16(Product2_acc_532_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_377_itm_17_2_1[15:1]) + conv_s2s_15_16(Product2_acc_127_cse_sva_1[15:1])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1)
      + conv_s2s_12_16(input_1_rsci_idat[79:68]) + 16'b1111111001000001;
  assign Product2_acc_1247_nl = nl_Product2_acc_1247_nl[15:0];
  assign nl_Product2_acc_1245_nl = (~ (input_1_rsci_idat[79:64])) + conv_s2s_15_16(Product2_acc_867_cse_sva_1[15:1]);
  assign Product2_acc_1245_nl = nl_Product2_acc_1245_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1 = Product2_acc_1248_nl
      + Product2_acc_1247_nl + Product2_acc_1245_nl + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_456_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_330_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[143:132]);
  assign Accum2_acc_330_nl = nl_Accum2_acc_330_nl[12:0];
  assign nl_Accum2_acc_1550_nl = conv_s2s_4_5(input_1_rsci_idat[223:220]) + 5'b00001;
  assign Accum2_acc_1550_nl = nl_Accum2_acc_1550_nl[4:0];
  assign nl_Accum2_acc_338_nl = conv_s2s_15_16(Product2_acc_667_cse_sva_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(Accum2_acc_330_nl) + conv_s2s_13_16({Accum2_acc_1550_nl ,
      (input_1_rsci_idat[219:212])});
  assign Accum2_acc_338_nl = nl_Accum2_acc_338_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1 = Accum2_acc_338_nl
      + conv_s2s_14_16(Product2_acc_447_itm_15_1_1[14:1]) + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_122_itm_17_2_1[15:2]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_347_nl = Product2_acc_937_itm_18_3_1 + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2])
      + conv_s2s_13_16(input_1_rsci_idat[95:83]) + conv_s2s_13_16(input_1_rsci_idat[175:163]);
  assign Accum2_acc_347_nl = nl_Accum2_acc_347_nl[15:0];
  assign nl_Accum2_acc_350_nl = Accum2_acc_347_nl + conv_s2s_15_16(Accum2_acc_343_cse_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_350_nl = nl_Accum2_acc_350_nl[15:0];
  assign nl_Accum2_acc_1551_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1[12:7])
      + 6'b111111;
  assign Accum2_acc_1551_nl = nl_Accum2_acc_1551_nl[5:0];
  assign nl_Accum2_acc_342_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1551_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1[6:0])});
  assign Accum2_acc_342_nl = nl_Accum2_acc_342_nl[13:0];
  assign nl_Accum2_acc_345_nl = conv_s2s_15_16(Product2_acc_1332_itm_17_2_1[15:1])
      + conv_s2s_14_16(Accum2_acc_342_nl);
  assign Accum2_acc_345_nl = nl_Accum2_acc_345_nl[15:0];
  assign nl_Product2_acc_1041_nl = conv_s2u_13_17(input_1_rsci_idat[47:35]) + conv_s2u_16_17(input_1_rsci_idat[47:32]);
  assign Product2_acc_1041_nl = nl_Product2_acc_1041_nl[16:0];
  assign nl_Accum2_acc_349_nl = Accum2_acc_345_nl + (readslicef_17_16_1(Product2_acc_1041_nl));
  assign Accum2_acc_349_nl = nl_Accum2_acc_349_nl[15:0];
  assign nl_Accum2_acc_348_nl = Product2_acc_283_itm_18_3_1 + Product2_acc_609_cse_sva_1;
  assign Accum2_acc_348_nl = nl_Accum2_acc_348_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1 = Accum2_acc_350_nl
      + Accum2_acc_349_nl + Accum2_acc_348_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[14:10]!=5'b00000);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_174_nl = conv_s2s_15_16(~
      (input_1_rsci_idat[175:161])) + conv_s2s_15_16(Product2_acc_1330_itm_17_3_1)
      + conv_s2s_15_16(Product2_acc_458_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_290_itm_15_1_1);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_174_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_174_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_168_nl = conv_s2s_15_16(Product2_acc_8_itm_18_3_1[15:1])
      + conv_s2s_14_16(Product2_acc_934_itm_17_2_1[15:2]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_168_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_168_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_173_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_168_nl
      + Product2_acc_204_cse_sva_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_173_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_173_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_166_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1
      + conv_s2s_10_13({9'b100000000 , (~ (input_1_rsci_idat[160]))});
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_166_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_166_nl[12:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_174_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_173_nl + Product2_acc_374_itm_19_4_1
      + Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(input_1_rsci_idat[143:129]) + conv_s2s_14_16(Product2_acc_122_itm_17_2_1[15:2])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_166_nl);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_361_nl = conv_s2s_15_16(Product2_acc_801_itm_18_4_1) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_122_itm_17_2_1[15:1]);
  assign Accum2_acc_361_nl = nl_Accum2_acc_361_nl[15:0];
  assign nl_Accum2_acc_1552_nl = conv_s2s_6_7(input_1_rsci_idat[175:170]) + 7'b1111111;
  assign Accum2_acc_1552_nl = nl_Accum2_acc_1552_nl[6:0];
  assign nl_Accum2_acc_353_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1552_nl , (input_1_rsci_idat[169:164])});
  assign Accum2_acc_353_nl = nl_Accum2_acc_353_nl[13:0];
  assign nl_Accum2_acc_360_nl = conv_s2s_15_16(Product2_acc_8_itm_18_3_1[15:1]) +
      conv_s2s_14_16(Accum2_acc_353_nl) + conv_s2s_14_16(input_1_rsci_idat[63:50])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_360_nl = nl_Accum2_acc_360_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1 = Accum2_acc_361_nl
      + Accum2_acc_360_nl + conv_s2s_15_16(input_1_rsci_idat[159:145]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[14:10]!=5'b00000);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_186_nl = conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1])
      + conv_s2s_15_16(input_1_rsci_idat[191:177]) + conv_s2s_15_16(Product2_acc_629_itm_17_3_1)
      + conv_s2s_15_16(Product2_acc_1064_itm_16_1_1[15:1]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_186_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_186_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_179_nl = conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_127_cse_sva_1[15:1]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_179_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_179_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_185_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_179_nl
      + (~ (input_1_rsci_idat[15:0]));
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_185_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_185_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_184_nl = Product2_acc_191_itm_19_4_1
      + Product2_acc_459_cse_sva_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_184_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_184_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_183_nl = Product2_acc_538_cse_sva_1
      + Product2_acc_670_itm_19_4_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_183_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_183_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_178_nl = conv_s2s_14_15(Product2_acc_730_cse_sva_1[15:2])
      + conv_s2s_12_15(input_1_rsci_idat[31:20]) + 15'b111111010000001;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_178_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_178_nl[14:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_182_nl = Product2_acc_942_itm_17_2_1
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_acc_178_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_182_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_182_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_186_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_185_nl + nnet_product_mult_input_t_config2_weight_t_product_acc_184_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_183_nl + nnet_product_mult_input_t_config2_weight_t_product_acc_182_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_372_nl = Accum2_acc_285_cse_1 + conv_s2s_15_16(Product2_acc_871_itm_17_2_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_372_nl = nl_Accum2_acc_372_nl[15:0];
  assign nl_Accum2_acc_364_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_119_12_6 , (input_1_rsci_idat[137:132])});
  assign Accum2_acc_364_nl = nl_Accum2_acc_364_nl[13:0];
  assign nl_Accum2_acc_371_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(Accum2_acc_364_nl) + conv_s2s_14_16(Product2_acc_943_cse_sva_1[15:2]);
  assign Accum2_acc_371_nl = nl_Accum2_acc_371_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1 = Accum2_acc_372_nl
      + Accum2_acc_371_nl + conv_s2s_14_16(Product2_acc_733_itm_17_2_1[15:2]) + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2])
      + conv_s2s_14_16(input_1_rsci_idat[159:146]) + conv_s2s_14_16(Product2_acc_377_itm_17_2_1[15:2]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1554_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1[12:9])
      + 4'b1111;
  assign Accum2_acc_1554_nl = nl_Accum2_acc_1554_nl[3:0];
  assign nl_Accum2_acc_384_nl = conv_s2s_15_16(Product2_acc_671_itm_18_3_1[15:1])
      + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2]) + conv_s2s_13_16({Accum2_acc_1554_nl
      , (nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1[8:0])})
      + conv_s2s_14_16(Product2_acc_730_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_603_itm_15_1_1[14:1])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_384_nl = nl_Accum2_acc_384_nl[15:0];
  assign nl_Accum2_acc_383_nl = Product2_acc_1066_itm_16_1_1 + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_383_nl = nl_Accum2_acc_383_nl[15:0];
  assign nl_Accum2_acc_379_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_15(input_1_rsci_idat[191:179]) + conv_s2s_13_15(input_1_rsci_idat[207:195]);
  assign Accum2_acc_379_nl = nl_Accum2_acc_379_nl[14:0];
  assign nl_Accum2_acc_382_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Accum2_acc_379_nl);
  assign Accum2_acc_382_nl = nl_Accum2_acc_382_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1 = Accum2_acc_384_nl
      + Accum2_acc_383_nl + Accum2_acc_382_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_390_nl = conv_s2s_15_16(input_1_rsci_idat[191:177]) + conv_s2s_14_16(input_1_rsci_idat[47:34])
      + conv_s2s_12_16(input_1_rsci_idat[143:132]) + conv_s2s_12_16(input_1_rsci_idat[207:196]);
  assign Accum2_acc_390_nl = nl_Accum2_acc_390_nl[15:0];
  assign nl_Accum2_acc_394_nl = Accum2_acc_390_nl + Product2_acc_11_itm_17_2_1;
  assign Accum2_acc_394_nl = nl_Accum2_acc_394_nl[15:0];
  assign nl_Accum2_acc_389_nl = (Product2_acc_379_itm_18_3_1[15:1]) + conv_s2s_14_15(Accum2_acc_387_cse_1);
  assign Accum2_acc_389_nl = nl_Accum2_acc_389_nl[14:0];
  assign nl_Accum2_acc_391_nl = Product2_acc_937_itm_18_3_1 + conv_s2s_15_16(Accum2_acc_389_nl);
  assign Accum2_acc_391_nl = nl_Accum2_acc_391_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1 = Accum2_acc_394_nl
      + Accum2_acc_391_nl + Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_541_itm_19_4_1 + Product2_acc_191_itm_19_4_1 + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1555_nl = conv_s2s_8_9(Product2_acc_532_cse_sva_1[15:8]) +
      9'b111111101;
  assign Accum2_acc_1555_nl = nl_Accum2_acc_1555_nl[8:0];
  assign nl_Accum2_acc_405_nl = conv_s2s_15_16({Accum2_acc_1555_nl , (Product2_acc_532_cse_sva_1[7:2])})
      + conv_s2s_15_16(Product2_acc_876_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_946_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_801_itm_18_4_1);
  assign Accum2_acc_405_nl = nl_Accum2_acc_405_nl[15:0];
  assign nl_Accum2_acc_404_nl = Accum2_acc_399_cse_1 + Product2_acc_124_cse_sva_1;
  assign Accum2_acc_404_nl = nl_Accum2_acc_404_nl[15:0];
  assign nl_Accum2_acc_403_nl = Product2_acc_1066_itm_16_1_1 + Product2_acc_367_itm_19_4_1;
  assign Accum2_acc_403_nl = nl_Accum2_acc_403_nl[15:0];
  assign nl_Accum2_acc_398_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_398_nl = nl_Accum2_acc_398_nl[14:0];
  assign nl_Accum2_acc_402_nl = Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Accum2_acc_398_nl);
  assign Accum2_acc_402_nl = nl_Accum2_acc_402_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1 = Accum2_acc_405_nl
      + Accum2_acc_404_nl + Accum2_acc_403_nl + Accum2_acc_402_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_415_nl = Product2_acc_281_itm_19_4_1 + Product2_acc_370_cse_sva_1;
  assign Accum2_acc_415_nl = nl_Accum2_acc_415_nl[15:0];
  assign nl_Accum2_acc_414_nl = Product2_acc_742_itm_17_2_1 + Product2_acc_1126_itm_16_1_1;
  assign Accum2_acc_414_nl = nl_Accum2_acc_414_nl[15:0];
  assign nl_Accum2_acc_418_nl = Accum2_acc_415_nl + Accum2_acc_414_nl;
  assign Accum2_acc_418_nl = nl_Accum2_acc_418_nl[15:0];
  assign nl_Accum2_acc_409_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1);
  assign Accum2_acc_409_nl = nl_Accum2_acc_409_nl[13:0];
  assign nl_Accum2_acc_1556_nl = conv_s2s_5_6(input_1_rsci_idat[127:123]) + 6'b111111;
  assign Accum2_acc_1556_nl = nl_Accum2_acc_1556_nl[5:0];
  assign nl_Accum2_acc_417_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(input_1_rsci_idat[15:1]) + conv_s2s_14_16(Accum2_acc_409_nl)
      + conv_s2s_14_16({Accum2_acc_1556_nl , (input_1_rsci_idat[122:115])});
  assign Accum2_acc_417_nl = nl_Accum2_acc_417_nl[15:0];
  assign nl_Accum2_acc_416_nl = Accum2_acc_411_cse_1 + Product2_acc_195_cse_sva_1;
  assign Accum2_acc_416_nl = nl_Accum2_acc_416_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1 = Accum2_acc_418_nl
      + Accum2_acc_417_nl + Accum2_acc_416_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_421_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1);
  assign Accum2_acc_421_nl = nl_Accum2_acc_421_nl[13:0];
  assign nl_Accum2_acc_428_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_943_cse_sva_1[15:1]) + conv_s2s_15_16(Product2_acc_382_cse_sva_1[15:1])
      + conv_s2s_14_16(Accum2_acc_421_nl);
  assign Accum2_acc_428_nl = nl_Accum2_acc_428_nl[15:0];
  assign nl_Accum2_acc_1557_nl = conv_s2s_7_8(input_1_rsci_idat[31:25]) + 8'b00000101;
  assign Accum2_acc_1557_nl = nl_Accum2_acc_1557_nl[7:0];
  assign nl_Accum2_acc_422_nl = conv_s2s_14_15({Accum2_acc_1557_nl , (input_1_rsci_idat[24:19])})
      + conv_s2s_14_15(Product2_acc_603_itm_15_1_1[14:1]);
  assign Accum2_acc_422_nl = nl_Accum2_acc_422_nl[14:0];
  assign nl_Accum2_acc_425_nl = Product2_acc_743_cse_sva_1 + conv_s2s_15_16(Accum2_acc_422_nl);
  assign Accum2_acc_425_nl = nl_Accum2_acc_425_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1 = Accum2_acc_428_nl
      + Accum2_acc_426_cse_1 + Accum2_acc_425_nl + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[14:10]!=5'b00000);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_59_nl = ~((input_1_rsci_idat[67:64]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_195_nl = (Product2_acc_212_itm_18_3_1[15:1])
      + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1)
      + conv_s2s_12_15(input_1_rsci_idat[175:164]) + conv_s2s_9_15({8'b10100000 ,
      nnet_product_mult_input_t_config2_weight_t_product_nor_59_nl});
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_195_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_195_nl[14:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_198_nl = Product2_acc_601_itm_19_4_1
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_acc_195_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_198_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_198_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_191_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1
      + conv_s2s_12_13(~ (input_1_rsci_idat[79:68]));
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_191_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_191_nl[12:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_201_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_198_nl
      + conv_s2s_14_16(input_1_rsci_idat[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_124_cse_sva_1[15:2]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_191_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_201_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_201_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_200_nl = Product2_acc_73_itm_19_4_1
      + conv_s2s_15_16(Product2_acc_937_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_1330_itm_17_3_1);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_200_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_200_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_199_nl = Product2_acc_458_itm_18_3_1
      + Product2_acc_1095_itm_16_1_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_199_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_199_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_201_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_200_nl + nnet_product_mult_input_t_config2_weight_t_product_acc_199_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_441_nl = conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1])
      + conv_s2s_15_16(Product2_acc_1095_itm_16_1_1[15:1]) + conv_s2s_14_16(Product2_acc_603_itm_15_1_1[14:1])
      + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_124_cse_sva_1[15:2])
      + conv_s2s_14_16(Product2_acc_297_itm_17_2_1[15:2]);
  assign Accum2_acc_441_nl = nl_Accum2_acc_441_nl[15:0];
  assign nl_Accum2_acc_440_nl = Product2_acc_450_itm_19_4_1 + conv_s2s_15_16(Product2_acc_1338_itm_17_3_1)
      + conv_s2s_13_16({Accum2_acc_1558_cse_1 , (input_1_rsci_idat[25:20])}) + conv_s2s_13_16(input_1_rsci_idat[159:147]);
  assign Accum2_acc_440_nl = nl_Accum2_acc_440_nl[15:0];
  assign nl_Accum2_acc_439_nl = Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_730_cse_sva_1[15:2]);
  assign Accum2_acc_439_nl = nl_Accum2_acc_439_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1 = Accum2_acc_441_nl
      + Accum2_acc_440_nl + Accum2_acc_439_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_446_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_12_14(input_1_rsci_idat[79:68]) + conv_s2s_12_14(input_1_rsci_idat[111:100]);
  assign Accum2_acc_446_nl = nl_Accum2_acc_446_nl[13:0];
  assign nl_Accum2_acc_1559_nl = conv_s2s_5_6(input_1_rsci_idat[127:123]) + 6'b111101;
  assign Accum2_acc_1559_nl = nl_Accum2_acc_1559_nl[5:0];
  assign nl_Accum2_acc_452_nl = Product2_acc_932_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_446_nl)
      + conv_s2s_13_16({Accum2_acc_1559_nl , (input_1_rsci_idat[122:116])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_452_nl = nl_Accum2_acc_452_nl[15:0];
  assign nl_Product2_acc_617_nl = conv_s2s_16_19(~ (input_1_rsci_idat[143:128]))
      + ({(input_1_rsci_idat[143:128]) , 3'b001});
  assign Product2_acc_617_nl = nl_Product2_acc_617_nl[18:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1 = Accum2_acc_452_nl
      + conv_s2s_15_16(Accum2_acc_447_cse_1) + conv_s2s_14_16(Product2_acc_1330_itm_17_3_1[14:1])
      + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(readslicef_19_15_4(Product2_acc_617_nl));
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1560_nl = conv_s2s_4_5(input_1_rsci_idat[191:188]) + 5'b00011;
  assign Accum2_acc_1560_nl = nl_Accum2_acc_1560_nl[4:0];
  assign nl_Accum2_acc_463_nl = conv_s2s_15_16(Accum2_acc_457_cse_1) + conv_s2s_15_16(input_1_rsci_idat[127:113])
      + conv_s2s_15_16(Product2_acc_867_cse_sva_1[15:1]) + conv_s2s_14_16(Product2_acc_1338_itm_17_3_1[14:1])
      + conv_s2s_13_16({Accum2_acc_1560_nl , (input_1_rsci_idat[187:180])});
  assign Accum2_acc_463_nl = nl_Accum2_acc_463_nl[15:0];
  assign nl_Accum2_acc_458_nl = conv_s2s_15_16(Product2_acc_204_cse_sva_1[15:1])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1);
  assign Accum2_acc_458_nl = nl_Accum2_acc_458_nl[15:0];
  assign nl_Accum2_acc_462_nl = Accum2_acc_458_nl + Product2_acc_298_itm_17_2_1;
  assign Accum2_acc_462_nl = nl_Accum2_acc_462_nl[15:0];
  assign nl_Accum2_acc_461_nl = Product2_acc_370_cse_sva_1 + Product2_acc_458_itm_18_3_1;
  assign Accum2_acc_461_nl = nl_Accum2_acc_461_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1 = Accum2_acc_463_nl
      + Accum2_acc_462_nl + Accum2_acc_461_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_473_nl = conv_s2s_15_16(input_1_rsci_idat[111:97]) + conv_s2s_15_16(input_1_rsci_idat[223:209])
      + conv_s2s_15_16(Product2_acc_1095_itm_16_1_1[15:1]) + conv_s2s_15_16(Product2_acc_1042_itm_16_1_1[15:1]);
  assign Accum2_acc_473_nl = nl_Accum2_acc_473_nl[15:0];
  assign nl_Accum2_acc_1561_nl = conv_s2s_6_7(input_1_rsci_idat[15:10]) + 7'b1111111;
  assign Accum2_acc_1561_nl = nl_Accum2_acc_1561_nl[6:0];
  assign nl_Accum2_acc_471_nl = Product2_acc_374_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_387_cse_1)
      + conv_s2s_13_16({Accum2_acc_1561_nl , (input_1_rsci_idat[9:4])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1);
  assign Accum2_acc_471_nl = nl_Accum2_acc_471_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1 = Accum2_acc_473_nl
      + Accum2_acc_471_nl + Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1562_nl = conv_s2s_6_7(input_1_rsci_idat[15:10]) + 7'b0000001;
  assign Accum2_acc_1562_nl = nl_Accum2_acc_1562_nl[6:0];
  assign nl_Accum2_acc_484_nl = conv_s2s_15_16(Product2_acc_667_cse_sva_1[15:1])
      + conv_s2s_13_16({Accum2_acc_1562_nl , (input_1_rsci_idat[9:4])}) + conv_s2s_13_16(input_1_rsci_idat[47:35])
      + conv_s2s_14_16(Accum2_acc_476_cse_1) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_603_itm_15_1_1[14:1]);
  assign Accum2_acc_484_nl = nl_Accum2_acc_484_nl[15:0];
  assign nl_Accum2_acc_483_nl = Product2_acc_214_cse_sva_1 + Product2_acc_429_itm_18_3_1;
  assign Accum2_acc_483_nl = nl_Accum2_acc_483_nl[15:0];
  assign nl_Accum2_acc_482_nl = Product2_acc_456_itm_19_4_1 + Product2_acc_547_itm_17_2_1;
  assign Accum2_acc_482_nl = nl_Accum2_acc_482_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1 = Accum2_acc_484_nl
      + Accum2_acc_483_nl + Accum2_acc_482_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_490_nl = Product2_acc_382_cse_sva_1 + Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_490_nl = nl_Accum2_acc_490_nl[15:0];
  assign nl_Accum2_acc_487_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[63:52]);
  assign Accum2_acc_487_nl = nl_Accum2_acc_487_nl[12:0];
  assign nl_Accum2_acc_1563_nl = conv_s2s_6_7(input_1_rsci_idat[223:218]) + 7'b1110101;
  assign Accum2_acc_1563_nl = nl_Accum2_acc_1563_nl[6:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1 = Accum2_acc_490_nl
      + Product2_acc_299_itm_19_4_1 + conv_s2s_15_16(Product2_acc_1338_itm_17_3_1)
      + conv_s2s_13_16(Accum2_acc_487_nl) + conv_s2s_13_16({Accum2_acc_1563_nl ,
      (input_1_rsci_idat[217:212])});
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_501_nl = conv_s2s_15_16(Product2_acc_604_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_127_cse_sva_1[15:1]) + conv_s2s_15_16(Product2_acc_1027_itm_16_2_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_501_nl = nl_Accum2_acc_501_nl[15:0];
  assign nl_Accum2_acc_498_nl = Product2_acc_727_itm_19_4_1 + Product2_acc_867_cse_sva_1;
  assign Accum2_acc_498_nl = nl_Accum2_acc_498_nl[15:0];
  assign nl_Accum2_acc_1564_nl = conv_s2s_6_7(input_1_rsci_idat[191:186]) + 7'b0000011;
  assign Accum2_acc_1564_nl = nl_Accum2_acc_1564_nl[6:0];
  assign nl_Accum2_acc_493_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1564_nl , (input_1_rsci_idat[185:180])});
  assign Accum2_acc_493_nl = nl_Accum2_acc_493_nl[13:0];
  assign nl_Accum2_acc_497_nl = Product2_acc_951_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_493_nl)
      + conv_s2s_14_16(Product2_acc_667_cse_sva_1[15:2]);
  assign Accum2_acc_497_nl = nl_Accum2_acc_497_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1 = Accum2_acc_501_nl
      + Accum2_acc_426_cse_1 + Product2_acc_212_itm_18_3_1 + Product2_acc_379_itm_18_3_1
      + Accum2_acc_498_nl + Accum2_acc_497_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[14:10]!=5'b00000);
  assign Product2_acc_1320_nl =  -conv_s2s_13_14(input_1_rsci_idat[159:147]);
  assign nl_Product2_acc_678_nl = conv_s2s_17_20({Product2_acc_1320_nl , (~ (input_1_rsci_idat[146:144]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[159:144])) , 3'b001});
  assign Product2_acc_678_nl = nl_Product2_acc_678_nl[19:0];
  assign nl_Accum2_acc_513_nl = Product2_acc_609_cse_sva_1 + (readslicef_20_16_4(Product2_acc_678_nl));
  assign Accum2_acc_513_nl = nl_Accum2_acc_513_nl[15:0];
  assign nl_Accum2_acc_512_nl = conv_s2s_15_16(Product2_acc_733_itm_17_2_1[15:1])
      + conv_s2s_14_16(Product2_acc_867_cse_sva_1[15:2]) + conv_s2s_13_16(input_1_rsci_idat[31:19])
      + conv_s2s_13_16(input_1_rsci_idat[79:67]);
  assign Accum2_acc_512_nl = nl_Accum2_acc_512_nl[15:0];
  assign nl_Accum2_acc_516_nl = Accum2_acc_513_nl + Accum2_acc_512_nl;
  assign Accum2_acc_516_nl = nl_Accum2_acc_516_nl[15:0];
  assign nl_Accum2_acc_1565_nl = conv_s2s_4_5(input_1_rsci_idat[223:220]) + 5'b00011;
  assign Accum2_acc_1565_nl = nl_Accum2_acc_1565_nl[4:0];
  assign nl_Accum2_acc_515_nl = conv_s2s_15_16(Product2_acc_1095_itm_16_1_1[15:1])
      + conv_s2s_15_16(Product2_acc_1079_itm_16_1_1[15:1]) + conv_s2s_15_16(Product2_acc_216_itm_18_3_1[15:1])
      + conv_s2s_13_16({Accum2_acc_1565_nl , (input_1_rsci_idat[219:212])}) + conv_s2s_12_16(input_1_rsci_idat[111:100])
      + conv_s2s_12_16(input_1_rsci_idat[191:180]);
  assign Accum2_acc_515_nl = nl_Accum2_acc_515_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1 = Accum2_acc_516_nl
      + Accum2_acc_515_nl + Product2_acc_itm_18_3_1 + Product2_acc_141_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_529_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_1110_itm_16_2_1) + conv_s2s_15_16(Product2_acc_532_cse_sva_1[15:1])
      + conv_s2s_14_16(Product2_acc_217_itm_17_2_1[15:2]) + conv_s2s_13_16(input_1_rsci_idat[31:19]);
  assign Accum2_acc_529_nl = nl_Accum2_acc_529_nl[15:0];
  assign nl_Accum2_acc_528_nl = conv_s2s_15_16(Product2_acc_1064_itm_16_1_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_3_itm_15_1_1) + conv_s2s_13_16(input_1_rsci_idat[143:131])
      + conv_s2s_13_16(input_1_rsci_idat[175:163]);
  assign Accum2_acc_528_nl = nl_Accum2_acc_528_nl[15:0];
  assign nl_Accum2_acc_1566_nl = conv_s2s_7_8(input_1_rsci_idat[223:217]) + 8'b00000001;
  assign Accum2_acc_1566_nl = nl_Accum2_acc_1566_nl[7:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1 = Accum2_acc_529_nl
      + Accum2_acc_528_nl + conv_s2s_14_16({Accum2_acc_1566_nl , (input_1_rsci_idat[216:211])})
      + conv_s2s_14_16(input_1_rsci_idat[111:98]) + conv_s2s_14_16(input_1_rsci_idat[191:178])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_536_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(Accum2_acc_532_cse_1);
  assign Accum2_acc_536_nl = nl_Accum2_acc_536_nl[13:0];
  assign nl_Accum2_acc_1567_nl = conv_s2s_6_7(input_1_rsci_idat[159:154]) + 7'b0001001;
  assign Accum2_acc_1567_nl = nl_Accum2_acc_1567_nl[6:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1 = Product2_acc_75_itm_19_4_1
      + Product2_acc_952_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_534_cse_1) + conv_s2s_14_16(input_1_rsci_idat[95:82])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_887_itm_15_1_1) + conv_s2s_14_16(Accum2_acc_536_nl)
      + conv_s2s_13_16({Accum2_acc_1567_nl , (input_1_rsci_idat[153:148])}) + conv_s2s_13_16(input_1_rsci_idat[47:35]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_552_nl = conv_s2s_15_16(Product2_acc_447_itm_15_1_1) + conv_s2s_15_16(Product2_acc_377_itm_17_2_1[15:1])
      + conv_s2s_13_16({Accum2_Accum2_conc_121_12_8 , (input_1_rsci_idat[219:212])})
      + conv_s2s_13_16(input_1_rsci_idat[79:67]) + conv_s2s_13_16(input_1_rsci_idat[127:115])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1);
  assign Accum2_acc_552_nl = nl_Accum2_acc_552_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1 = Accum2_acc_552_nl
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_217_itm_17_2_1[15:2]) + conv_s2s_14_16(Product2_acc_1338_itm_17_3_1[14:1]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[14:10]!=5'b00000);
  assign Product2_acc_1321_nl =  -conv_s2s_12_13(input_1_rsci_idat[175:164]);
  assign nl_Product2_acc_1253_nl = ({(input_1_rsci_idat[175:160]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1321_nl
      , (~ (input_1_rsci_idat[163:160]))});
  assign Product2_acc_1253_nl = nl_Product2_acc_1253_nl[17:0];
  assign nl_Product2_acc_747_nl = conv_s2s_18_20(Product2_acc_1253_nl) + ({(~ (input_1_rsci_idat[175:160]))
      , 4'b0000});
  assign Product2_acc_747_nl = nl_Product2_acc_747_nl[19:0];
  assign nl_Accum2_acc_559_nl = Product2_acc_458_itm_18_3_1 + (readslicef_20_16_4(Product2_acc_747_nl));
  assign Accum2_acc_559_nl = nl_Accum2_acc_559_nl[15:0];
  assign nl_Product2_acc_1254_nl = (~ (input_1_rsci_idat[223:208])) + conv_s2s_14_16(input_1_rsci_idat[223:210]);
  assign Product2_acc_1254_nl = nl_Product2_acc_1254_nl[15:0];
  assign nl_Product2_acc_1146_nl = conv_s2u_16_18(Product2_acc_1254_nl) + ({(input_1_rsci_idat[223:208])
      , 2'b01});
  assign Product2_acc_1146_nl = nl_Product2_acc_1146_nl[17:0];
  assign nl_Accum2_acc_558_nl = Product2_acc_1126_itm_16_1_1 + (readslicef_18_16_2(Product2_acc_1146_nl));
  assign Accum2_acc_558_nl = nl_Accum2_acc_558_nl[15:0];
  assign nl_Accum2_acc_562_nl = Accum2_acc_559_nl + Accum2_acc_558_nl;
  assign Accum2_acc_562_nl = nl_Accum2_acc_562_nl[15:0];
  assign nl_Accum2_acc_555_nl = (Product2_acc_379_itm_18_3_1[15:1]) + conv_s2s_13_15(input_1_rsci_idat[143:131])
      + conv_s2s_12_15(input_1_rsci_idat[207:196]);
  assign Accum2_acc_555_nl = nl_Accum2_acc_555_nl[14:0];
  assign nl_Accum2_acc_561_nl = conv_s2s_15_16(Accum2_acc_555_nl) + conv_s2s_15_16(Product2_acc_1330_itm_17_3_1)
      + conv_s2s_15_16(Product2_acc_1095_itm_16_1_1[15:1]) + conv_s2s_14_16(Product2_acc_1338_itm_17_3_1[14:1])
      + conv_s2s_13_16(input_1_rsci_idat[31:19]);
  assign Accum2_acc_561_nl = nl_Accum2_acc_561_nl[15:0];
  assign nl_Accum2_acc_560_nl = Product2_acc_141_itm_19_4_1 + Product2_acc_1053_itm_16_1_1;
  assign Accum2_acc_560_nl = nl_Accum2_acc_560_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1 = Accum2_acc_562_nl
      + Accum2_acc_561_nl + Accum2_acc_560_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1569_nl = conv_s2s_5_6(input_1_rsci_idat[15:11]) + 6'b000001;
  assign Accum2_acc_1569_nl = nl_Accum2_acc_1569_nl[5:0];
  assign nl_Accum2_acc_568_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_15({Accum2_acc_1569_nl , (input_1_rsci_idat[10:4])}) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1);
  assign Accum2_acc_568_nl = nl_Accum2_acc_568_nl[14:0];
  assign nl_Accum2_acc_574_nl = conv_s2s_15_16(Accum2_acc_568_nl) + conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_447_itm_15_1_1[14:1]) + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_574_nl = nl_Accum2_acc_574_nl[15:0];
  assign nl_Accum2_acc_573_nl = Product2_acc_1336_itm_18_3_1 + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_538_cse_sva_1[15:1]);
  assign Accum2_acc_573_nl = nl_Accum2_acc_573_nl[15:0];
  assign nl_Product2_acc_1104_nl = conv_s2u_13_17(input_1_rsci_idat[143:131]) + conv_s2u_16_17(input_1_rsci_idat[143:128]);
  assign Product2_acc_1104_nl = nl_Product2_acc_1104_nl[16:0];
  assign nl_Accum2_acc_572_nl = (readslicef_17_16_1(Product2_acc_1104_nl)) + Product2_acc_954_itm_19_4_1;
  assign Accum2_acc_572_nl = nl_Accum2_acc_572_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1 = Accum2_acc_574_nl
      + Accum2_acc_573_nl + Accum2_acc_572_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_585_nl = Product2_acc_191_itm_19_4_1 + conv_s2s_15_16(input_1_rsci_idat[175:161])
      + conv_s2s_15_16(Product2_acc_532_cse_sva_1[15:1]);
  assign Accum2_acc_585_nl = nl_Accum2_acc_585_nl[15:0];
  assign nl_Accum2_acc_584_nl = Product2_acc_281_itm_19_4_1 + Product2_acc_394_itm_17_2_1;
  assign Accum2_acc_584_nl = nl_Accum2_acc_584_nl[15:0];
  assign nl_Accum2_acc_1570_nl = conv_s2s_3_4(input_1_rsci_idat[111:109]) + 4'b0001;
  assign Accum2_acc_1570_nl = nl_Accum2_acc_1570_nl[3:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1 = Accum2_acc_585_nl
      + Accum2_acc_584_nl + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_809_itm_19_4_1 + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_1338_itm_17_3_1[14:1]) + conv_s2s_13_16({Accum2_acc_1570_nl
      , (input_1_rsci_idat[108:100])}) + conv_s2s_13_16(input_1_rsci_idat[159:147])
      + conv_s2s_13_16(input_1_rsci_idat[207:195]) + conv_s2s_12_16(input_1_rsci_idat[47:36]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_595_nl = Accum2_acc_590_cse_1 + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_1086_itm_16_1_1[15:1]);
  assign Accum2_acc_595_nl = nl_Accum2_acc_595_nl[15:0];
  assign nl_Accum2_acc_594_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_1064_itm_16_1_1;
  assign Accum2_acc_594_nl = nl_Accum2_acc_594_nl[15:0];
  assign nl_Accum2_acc_1571_nl = (Product2_acc_1338_itm_17_3_1[14:7]) + 8'b11111111;
  assign Accum2_acc_1571_nl = nl_Accum2_acc_1571_nl[7:0];
  assign nl_Accum2_acc_589_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15({Accum2_acc_1571_nl , (Product2_acc_1338_itm_17_3_1[6:1])});
  assign Accum2_acc_589_nl = nl_Accum2_acc_589_nl[14:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1 = Accum2_acc_595_nl
      + Accum2_acc_594_nl + Product2_acc_606_itm_19_4_1 + Product2_acc_952_itm_19_4_1
      + conv_s2s_15_16(Accum2_acc_589_nl) + conv_s2s_15_16(Product2_acc_666_itm_18_3_1[15:1]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[14:10]!=5'b00000);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_213_nl = conv_s2s_15_16(~
      (input_1_rsci_idat[191:177])) + conv_s2s_15_16(Product2_acc_1330_itm_17_3_1)
      + conv_s2s_15_16(Product2_acc_283_itm_18_3_1[15:1]) + conv_s2s_14_16(Product2_acc_733_itm_17_2_1[15:2])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_213_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_213_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_212_nl = Product2_acc_217_itm_17_2_1
      + conv_s2s_15_16(Product2_acc_379_itm_18_3_1[15:1]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_212_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_212_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_210_nl = Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1)
      + conv_s2s_12_16(input_1_rsci_idat[15:4]) + conv_s2s_9_16({8'b10000000 , (~
      (input_1_rsci_idat[176]))});
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_210_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_210_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_213_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_212_nl + nnet_product_mult_input_t_config2_weight_t_product_acc_210_nl
      + Product2_acc_450_itm_19_4_1 + Product2_acc_554_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_600_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[47:36]);
  assign Accum2_acc_600_nl = nl_Accum2_acc_600_nl[12:0];
  assign nl_Accum2_acc_603_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(Accum2_acc_600_nl);
  assign Accum2_acc_603_nl = nl_Accum2_acc_603_nl[13:0];
  assign nl_Accum2_acc_609_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_603_itm_15_1_1) + conv_s2s_15_16(Product2_acc_1086_itm_16_1_1[15:1])
      + conv_s2s_14_16(Accum2_acc_603_nl);
  assign Accum2_acc_609_nl = nl_Accum2_acc_609_nl[15:0];
  assign nl_Accum2_acc_1572_nl = conv_s2s_6_7(input_1_rsci_idat[159:154]) + 7'b0000001;
  assign Accum2_acc_1572_nl = nl_Accum2_acc_1572_nl[6:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1 = Accum2_acc_609_nl
      + Product2_acc_73_itm_19_4_1 + Product2_acc_531_itm_19_4_1 + conv_s2s_15_16(Product2_acc_887_itm_15_1_1)
      + conv_s2s_13_16({Accum2_acc_1572_nl , (input_1_rsci_idat[153:148])}) + conv_s2s_12_16(input_1_rsci_idat[63:52])
      + conv_s2s_12_16(input_1_rsci_idat[95:84]) + conv_s2s_13_16(input_1_rsci_idat[79:67])
      + conv_s2s_13_16(input_1_rsci_idat[175:163]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[14:10]!=5'b00000);
  assign Product2_acc_1322_nl =  -conv_s2s_12_13(input_1_rsci_idat[31:20]);
  assign nl_Product2_acc_1256_nl = ({(input_1_rsci_idat[31:16]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1322_nl
      , (~ (input_1_rsci_idat[19:16]))});
  assign Product2_acc_1256_nl = nl_Product2_acc_1256_nl[17:0];
  assign nl_Product2_acc_78_nl = conv_s2s_18_20(Product2_acc_1256_nl) + ({(~ (input_1_rsci_idat[31:16]))
      , 4'b0000});
  assign Product2_acc_78_nl = nl_Product2_acc_78_nl[19:0];
  assign nl_Accum2_acc_619_nl = (readslicef_20_16_4(Product2_acc_78_nl)) + Product2_acc_195_cse_sva_1;
  assign Accum2_acc_619_nl = nl_Accum2_acc_619_nl[15:0];
  assign nl_Accum2_acc_618_nl = Product2_acc_281_itm_19_4_1 + Product2_acc_367_itm_19_4_1;
  assign Accum2_acc_618_nl = nl_Accum2_acc_618_nl[15:0];
  assign nl_Accum2_acc_622_nl = Accum2_acc_619_nl + Accum2_acc_618_nl;
  assign Accum2_acc_622_nl = nl_Accum2_acc_622_nl[15:0];
  assign nl_Accum2_acc_620_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_743_cse_sva_1[15:1]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_620_nl = nl_Accum2_acc_620_nl[15:0];
  assign nl_Product2_acc_1257_nl = (~ (input_1_rsci_idat[159:144])) + conv_s2s_14_16(input_1_rsci_idat[159:146]);
  assign Product2_acc_1257_nl = nl_Product2_acc_1257_nl[15:0];
  assign nl_Product2_acc_1111_nl = conv_s2u_16_18(Product2_acc_1257_nl) + ({(input_1_rsci_idat[159:144])
      , 2'b01});
  assign Product2_acc_1111_nl = nl_Product2_acc_1111_nl[17:0];
  assign nl_Accum2_acc_617_nl = Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + (readslicef_18_16_2(Product2_acc_1111_nl));
  assign Accum2_acc_617_nl = nl_Accum2_acc_617_nl[15:0];
  assign nl_Accum2_acc_1573_nl = conv_s2s_4_5(input_1_rsci_idat[47:44]) + 5'b00001;
  assign Accum2_acc_1573_nl = nl_Accum2_acc_1573_nl[4:0];
  assign nl_Accum2_acc_612_nl = ({Accum2_acc_1573_nl , (input_1_rsci_idat[43:35])})
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1);
  assign Accum2_acc_612_nl = nl_Accum2_acc_612_nl[13:0];
  assign nl_Accum2_acc_613_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15(Accum2_acc_612_nl);
  assign Accum2_acc_613_nl = nl_Accum2_acc_613_nl[14:0];
  assign nl_Accum2_acc_616_nl = Product2_acc_943_cse_sva_1 + conv_s2s_15_16(Accum2_acc_613_nl);
  assign Accum2_acc_616_nl = nl_Accum2_acc_616_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1 = Accum2_acc_622_nl
      + Accum2_acc_620_nl + Accum2_acc_617_nl + Accum2_acc_616_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1574_nl = conv_s2s_6_7(input_1_rsci_idat[143:138]) + 7'b1111101;
  assign Accum2_acc_1574_nl = nl_Accum2_acc_1574_nl[6:0];
  assign nl_Accum2_acc_626_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1574_nl , (input_1_rsci_idat[137:132])});
  assign Accum2_acc_626_nl = nl_Accum2_acc_626_nl[13:0];
  assign nl_Accum2_acc_633_nl = conv_s2s_15_16(Product2_acc_1086_itm_16_1_1[15:1])
      + conv_s2s_14_16(Accum2_acc_626_nl) + conv_s2s_13_16(input_1_rsci_idat[63:51])
      + conv_s2s_13_16(input_1_rsci_idat[223:211]) + conv_s2s_14_16(input_1_rsci_idat[207:194])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_633_nl = nl_Accum2_acc_633_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1 = Accum2_acc_633_nl
      + conv_s2s_14_16(input_1_rsci_idat[47:34]) + conv_s2s_14_16(input_1_rsci_idat[79:66])
      + conv_s2s_14_16(input_1_rsci_idat[95:82]) + conv_s2s_14_16(input_1_rsci_idat[127:114]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_642_nl = Product2_acc_1056_itm_16_1_1 + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_642_nl = nl_Accum2_acc_642_nl[15:0];
  assign nl_Accum2_acc_637_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_113_12_9 , (input_1_rsci_idat[12:4])});
  assign Accum2_acc_637_nl = nl_Accum2_acc_637_nl[13:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1 = Accum2_acc_642_nl
      + Product2_acc_398_itm_19_4_1 + Product2_acc_478_itm_17_2_1 + conv_s2s_14_16(Accum2_acc_637_nl)
      + conv_s2s_14_16(Accum2_acc_635_cse_1) + conv_s2s_14_16(Product2_acc_934_itm_17_2_1[15:2])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[14:10]!=5'b00000);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_223_nl = Product2_acc_1114_itm_17_2_1
      + Product2_acc_1134_itm_16_1_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_223_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_223_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_217_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[15:4]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_217_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_217_nl[12:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_219_nl = conv_s2s_14_15(Product2_acc_1330_itm_17_3_1[14:1])
      + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_217_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_219_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_219_nl[14:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_222_nl = Product2_acc_936_cse_sva_1
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_acc_219_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_222_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_222_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_226_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_223_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_222_nl;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_226_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_226_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_225_nl = conv_s2s_15_16(Product2_acc_532_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_603_itm_15_1_1) + conv_s2s_15_16(Product2_acc_308_cse_sva_1[15:1])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1)
      + conv_s2s_12_16(input_1_rsci_idat[47:36]) + 16'b1111111010000001;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_225_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_225_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_224_nl = (~ (input_1_rsci_idat[191:176]))
      + Product2_acc_191_itm_19_4_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_224_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_224_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_226_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_225_nl + nnet_product_mult_input_t_config2_weight_t_product_acc_224_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_652_nl = conv_s2s_15_16(input_1_rsci_idat[175:161]) + conv_s2s_15_16(Product2_acc_1105_itm_16_1_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_652_nl = nl_Accum2_acc_652_nl[15:0];
  assign nl_Accum2_acc_650_nl = Product2_acc_476_itm_19_4_1 + Product2_acc_1101_itm_16_1_1;
  assign Accum2_acc_650_nl = nl_Accum2_acc_650_nl[15:0];
  assign nl_Accum2_acc_1576_nl = conv_s2s_7_8(input_1_rsci_idat[207:201]) + 8'b11111011;
  assign Accum2_acc_1576_nl = nl_Accum2_acc_1576_nl[7:0];
  assign nl_Accum2_acc_649_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16({Accum2_acc_1576_nl , (input_1_rsci_idat[200:195])}) + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2]);
  assign Accum2_acc_649_nl = nl_Accum2_acc_649_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1 = Accum2_acc_652_nl
      + Accum2_acc_650_nl + Accum2_acc_649_nl + Product2_acc_212_itm_18_3_1 + Product2_acc_398_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_665_nl = conv_s2s_15_16(input_1_rsci_idat[79:65]) + conv_s2s_15_16(Product2_acc_665_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_379_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_itm_18_3_1[15:1]);
  assign Accum2_acc_665_nl = nl_Accum2_acc_665_nl[15:0];
  assign nl_Accum2_acc_664_nl = Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_216_itm_18_3_1[15:1]) + conv_s2s_13_16({Accum2_Accum2_conc_111_12_7
      , (input_1_rsci_idat[186:180])}) + conv_s2s_12_16(input_1_rsci_idat[47:36])
      + conv_s2s_12_16(input_1_rsci_idat[143:132]);
  assign Accum2_acc_664_nl = nl_Accum2_acc_664_nl[15:0];
  assign nl_Accum2_acc_663_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(input_1_rsci_idat[223:210]) + conv_s2s_13_16(input_1_rsci_idat[175:163])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_663_nl = nl_Accum2_acc_663_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1 = Accum2_acc_665_nl
      + Accum2_acc_664_nl + Accum2_acc_663_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1578_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1[12:8])
      + 5'b11111;
  assign Accum2_acc_1578_nl = nl_Accum2_acc_1578_nl[4:0];
  assign nl_Accum2_acc_669_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1578_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1[7:0])});
  assign Accum2_acc_669_nl = nl_Accum2_acc_669_nl[13:0];
  assign nl_Accum2_acc_671_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15(Accum2_acc_669_nl);
  assign Accum2_acc_671_nl = nl_Accum2_acc_671_nl[14:0];
  assign nl_Accum2_acc_673_nl = Product2_acc_932_itm_19_4_1 + conv_s2s_15_16(Accum2_acc_671_nl);
  assign Accum2_acc_673_nl = nl_Accum2_acc_673_nl[15:0];
  assign nl_Accum2_acc_676_nl = Accum2_acc_673_nl + conv_s2s_15_16(Product2_acc_665_cse_sva_1[15:1])
      + conv_s2s_14_16(input_1_rsci_idat[175:162]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1);
  assign Accum2_acc_676_nl = nl_Accum2_acc_676_nl[15:0];
  assign nl_Accum2_acc_674_nl = Product2_acc_367_itm_19_4_1 + Product2_acc_459_cse_sva_1;
  assign Accum2_acc_674_nl = nl_Accum2_acc_674_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1 = Accum2_acc_676_nl
      + Accum2_acc_674_nl + Product2_acc_212_itm_18_3_1 + Product2_acc_285_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_686_nl = Product2_acc_368_cse_sva_1 + Product2_acc_1134_itm_16_1_1;
  assign Accum2_acc_686_nl = nl_Accum2_acc_686_nl[15:0];
  assign nl_Accum2_acc_681_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15(Product2_acc_629_itm_17_3_1[14:1]);
  assign Accum2_acc_681_nl = nl_Accum2_acc_681_nl[14:0];
  assign nl_Accum2_acc_685_nl = conv_s2s_15_16(Accum2_acc_681_nl) + conv_s2s_14_16(Product2_acc_478_itm_17_2_1[15:2])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_685_nl = nl_Accum2_acc_685_nl[15:0];
  assign nl_Accum2_acc_689_nl = Accum2_acc_686_nl + Accum2_acc_685_nl;
  assign Accum2_acc_689_nl = nl_Accum2_acc_689_nl[15:0];
  assign nl_Accum2_acc_1579_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1[12:7])
      + 6'b111101;
  assign Accum2_acc_1579_nl = nl_Accum2_acc_1579_nl[5:0];
  assign nl_Accum2_acc_688_nl = conv_s2s_15_16(Product2_acc_1147_itm_16_2_1) + conv_s2s_15_16(Product2_acc_743_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_792_cse_sva_1[15:1]) + conv_s2s_14_16(Product2_acc_1332_itm_17_2_1[15:2])
      + conv_s2s_13_16({Accum2_acc_1579_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1[6:0])});
  assign Accum2_acc_688_nl = nl_Accum2_acc_688_nl[15:0];
  assign nl_Accum2_acc_687_nl = Product2_acc_141_itm_19_4_1 + conv_s2s_15_16(Product2_acc_308_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_217_itm_17_2_1[15:1]);
  assign Accum2_acc_687_nl = nl_Accum2_acc_687_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1 = Accum2_acc_689_nl
      + Accum2_acc_688_nl + Accum2_acc_687_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1580_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1[12:7])
      + 6'b000011;
  assign Accum2_acc_1580_nl = nl_Accum2_acc_1580_nl[5:0];
  assign nl_Accum2_acc_696_nl = Product2_acc_876_itm_18_3_1 + conv_s2s_14_16(input_1_rsci_idat[159:146])
      + conv_s2s_13_16({Accum2_acc_1580_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1[6:0])});
  assign Accum2_acc_696_nl = nl_Accum2_acc_696_nl[15:0];
  assign nl_Accum2_acc_700_nl = Accum2_acc_696_nl + conv_s2s_15_16(Product2_acc_934_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_447_itm_15_1_1);
  assign Accum2_acc_700_nl = nl_Accum2_acc_700_nl[15:0];
  assign nl_Accum2_acc_699_nl = conv_s2s_15_16(Product2_acc_560_itm_18_3_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_124_cse_sva_1[15:1]) + conv_s2s_14_16(input_1_rsci_idat[95:82]);
  assign Accum2_acc_699_nl = nl_Accum2_acc_699_nl[15:0];
  assign nl_Accum2_acc_697_nl = Product2_acc_1056_itm_16_1_1 + Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_697_nl = nl_Accum2_acc_697_nl[15:0];
  assign Product2_acc_1323_nl =  -conv_s2s_13_14(input_1_rsci_idat[15:3]);
  assign nl_Product2_acc_28_nl = conv_s2s_17_20({Product2_acc_1323_nl , (~ (input_1_rsci_idat[2:0]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[15:0])) , 3'b001});
  assign Product2_acc_28_nl = nl_Product2_acc_28_nl[19:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1 = Accum2_acc_700_nl
      + Accum2_acc_699_nl + Accum2_acc_697_nl + (readslicef_20_16_4(Product2_acc_28_nl))
      + Product2_acc_1332_itm_17_2_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[14:10]!=5'b00000);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_236_nl = Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(~ (input_1_rsci_idat[159:145])) + conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_236_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_236_nl[15:0];
  assign nl_Product2_acc_1259_nl = (~ (input_1_rsci_idat[143:128])) + conv_s2s_14_16(input_1_rsci_idat[143:130]);
  assign Product2_acc_1259_nl = nl_Product2_acc_1259_nl[15:0];
  assign nl_Product2_acc_1106_nl = conv_s2u_16_18(Product2_acc_1259_nl) + ({(input_1_rsci_idat[143:128])
      , 2'b01});
  assign Product2_acc_1106_nl = nl_Product2_acc_1106_nl[17:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_235_nl = Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + (readslicef_18_16_2(Product2_acc_1106_nl));
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_235_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_235_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_230_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_12_14(input_1_rsci_idat[63:52]) + conv_s2s_10_14({9'b101100000 ,
      (~ (input_1_rsci_idat[144]))});
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_230_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_230_nl[13:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_236_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_235_nl + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_acc_230_nl)
      + conv_s2s_14_16(Product2_acc_943_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_478_itm_17_2_1[15:2])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1581_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1[12:9])
      + 4'b1111;
  assign Accum2_acc_1581_nl = nl_Accum2_acc_1581_nl[3:0];
  assign nl_Accum2_acc_713_nl = conv_s2s_15_16(Product2_acc_478_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_290_itm_15_1_1) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_532_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_377_itm_17_2_1[15:2])
      + conv_s2s_13_16({Accum2_acc_1581_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1[8:0])});
  assign Accum2_acc_713_nl = nl_Accum2_acc_713_nl[15:0];
  assign nl_Accum2_acc_708_nl = conv_s2s_15_16(Product2_acc_1034_itm_16_1_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_708_nl = nl_Accum2_acc_708_nl[15:0];
  assign nl_Accum2_acc_712_nl = Accum2_acc_708_nl + Product2_acc_195_cse_sva_1;
  assign Accum2_acc_712_nl = nl_Accum2_acc_712_nl[15:0];
  assign nl_Accum2_acc_711_nl = Product2_acc_937_itm_18_3_1 + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2])
      + conv_s2s_13_16(input_1_rsci_idat[175:163]) + conv_s2s_13_16(input_1_rsci_idat[207:195]);
  assign Accum2_acc_711_nl = nl_Accum2_acc_711_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1 = Accum2_acc_713_nl
      + Accum2_acc_712_nl + Accum2_acc_711_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_724_nl = conv_s2s_15_16(Product2_acc_1126_itm_16_1_1[15:1])
      + conv_s2s_14_16(Product2_acc_85_itm_15_1_1[14:1]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[143:130]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_1338_itm_17_3_1[14:1]);
  assign Accum2_acc_724_nl = nl_Accum2_acc_724_nl[15:0];
  assign nl_Accum2_acc_1582_nl = conv_s2s_4_5(input_1_rsci_idat[79:76]) + 5'b00001;
  assign Accum2_acc_1582_nl = nl_Accum2_acc_1582_nl[4:0];
  assign nl_Accum2_acc_719_nl = (Product2_acc_379_itm_18_3_1[15:1]) + conv_s2s_14_15({Accum2_acc_1582_nl
      , (input_1_rsci_idat[75:67])});
  assign Accum2_acc_719_nl = nl_Accum2_acc_719_nl[14:0];
  assign nl_Accum2_acc_722_nl = Product2_acc_952_itm_19_4_1 + conv_s2s_15_16(Accum2_acc_719_nl);
  assign Accum2_acc_722_nl = nl_Accum2_acc_722_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1 = Accum2_acc_724_nl
      + Accum2_acc_722_nl + Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_734_nl = conv_s2s_15_16(input_1_rsci_idat[47:33]) + conv_s2s_15_16(Product2_acc_560_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_204_cse_sva_1[15:1]) + conv_s2s_14_16(Accum2_acc_727_cse_1);
  assign Accum2_acc_734_nl = nl_Accum2_acc_734_nl[15:0];
  assign nl_Accum2_acc_733_nl = Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[111:98]);
  assign Accum2_acc_733_nl = nl_Accum2_acc_733_nl[15:0];
  assign nl_Accum2_acc_1583_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[12:7])
      + 6'b111101;
  assign Accum2_acc_1583_nl = nl_Accum2_acc_1583_nl[5:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1 = Accum2_acc_734_nl
      + Accum2_acc_733_nl + conv_s2s_15_16(Product2_acc_1147_itm_16_2_1) + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2])
      + conv_s2s_13_16({Accum2_acc_1583_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[6:0])});
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[14:10]!=5'b00000);
  assign nl_Product2_acc_1264_nl = conv_s2s_14_15(input_1_rsci_idat[191:178]) + conv_s2s_14_15(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Product2_acc_1264_nl = nl_Product2_acc_1264_nl[14:0];
  assign nl_Product2_acc_1267_nl = (~ (input_1_rsci_idat[143:128])) + conv_s2s_15_16(Product2_acc_1264_nl);
  assign Product2_acc_1267_nl = nl_Product2_acc_1267_nl[15:0];
  assign nl_Product2_acc_1270_nl = Product2_acc_1267_nl + conv_s2s_15_16(Product2_acc_946_itm_18_3_1[15:1])
      + conv_s2s_14_16(Product2_acc_478_itm_17_2_1[15:2]) + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2]);
  assign Product2_acc_1270_nl = nl_Product2_acc_1270_nl[15:0];
  assign nl_Product2_acc_1261_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[95:84]);
  assign Product2_acc_1261_nl = nl_Product2_acc_1261_nl[12:0];
  assign nl_Product2_acc_1260_nl = conv_s2s_12_13(input_1_rsci_idat[143:132]) + 13'b0001001000001;
  assign Product2_acc_1260_nl = nl_Product2_acc_1260_nl[12:0];
  assign nl_Product2_acc_1265_nl = conv_s2s_15_16(Product2_acc_1064_itm_16_1_1[15:1])
      + conv_s2s_13_16(Product2_acc_1261_nl) + conv_s2s_13_16(Product2_acc_1260_nl);
  assign Product2_acc_1265_nl = nl_Product2_acc_1265_nl[15:0];
  assign nl_Product2_acc_1035_nl = conv_s2u_13_17(input_1_rsci_idat[31:19]) + conv_s2u_16_17(input_1_rsci_idat[31:16]);
  assign Product2_acc_1035_nl = nl_Product2_acc_1035_nl[16:0];
  assign nl_Product2_acc_1269_nl = Product2_acc_1265_nl + (readslicef_17_16_1(Product2_acc_1035_nl));
  assign Product2_acc_1269_nl = nl_Product2_acc_1269_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1 = Product2_acc_1270_nl
      + Product2_acc_1269_nl + Product2_acc_141_itm_19_4_1 + Product2_acc_691_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_746_nl = conv_s2s_15_16(Product2_acc_871_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_665_cse_sva_1[15:1]) + conv_s2s_13_16({Accum2_Accum2_conc_129_12_8
      , (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[7:0])})
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[127:115]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_308_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2]);
  assign Accum2_acc_746_nl = nl_Accum2_acc_746_nl[15:0];
  assign nl_Accum2_acc_741_nl = conv_s2s_15_16(Product2_acc_970_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_448_itm_15_1_1);
  assign Accum2_acc_741_nl = nl_Accum2_acc_741_nl[15:0];
  assign nl_Accum2_acc_745_nl = Accum2_acc_741_nl + Product2_acc_1042_itm_16_1_1;
  assign Accum2_acc_745_nl = nl_Accum2_acc_745_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1 = Accum2_acc_746_nl
      + Accum2_acc_745_nl + Product2_acc_193_itm_19_4_1 + Product2_acc_601_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_749_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[63:52]);
  assign Accum2_acc_749_nl = nl_Accum2_acc_749_nl[12:0];
  assign nl_Accum2_acc_1585_nl = conv_s2s_3_4(input_1_rsci_idat[223:221]) + 4'b1111;
  assign Accum2_acc_1585_nl = nl_Accum2_acc_1585_nl[3:0];
  assign nl_Accum2_acc_757_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(Product2_acc_730_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_1330_itm_17_3_1[14:1])
      + conv_s2s_13_16(Accum2_acc_749_nl) + conv_s2s_13_16({Accum2_acc_1585_nl ,
      (input_1_rsci_idat[220:212])});
  assign Accum2_acc_757_nl = nl_Accum2_acc_757_nl[15:0];
  assign nl_Accum2_acc_753_nl = conv_s2s_14_15(Product2_acc_867_cse_sva_1[15:2])
      + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1)
      + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1);
  assign Accum2_acc_753_nl = nl_Accum2_acc_753_nl[14:0];
  assign nl_Accum2_acc_755_nl = Product2_acc_1126_itm_16_1_1 + conv_s2s_15_16(Accum2_acc_753_nl);
  assign Accum2_acc_755_nl = nl_Accum2_acc_755_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1 = Accum2_acc_757_nl
      + Accum2_acc_755_nl + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[14:10]!=5'b00000);
  assign nl_Product2_acc_900_nl = conv_s2s_16_20(~ (input_1_rsci_idat[207:192]))
      + ({(input_1_rsci_idat[207:192]) , 4'b0001});
  assign Product2_acc_900_nl = nl_Product2_acc_900_nl[19:0];
  assign nl_Accum2_acc_769_nl = (readslicef_20_16_4(Product2_acc_900_nl)) + Product2_acc_954_itm_19_4_1
      + conv_s2s_14_16(Product2_acc_730_cse_sva_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[95:82]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_769_nl = nl_Accum2_acc_769_nl[15:0];
  assign nl_Accum2_acc_1586_nl = conv_s2s_4_5(input_1_rsci_idat[127:124]) + 5'b00001;
  assign Accum2_acc_1586_nl = nl_Accum2_acc_1586_nl[4:0];
  assign nl_Accum2_acc_768_nl = Product2_acc_1332_itm_17_2_1 + conv_s2s_15_16(Product2_acc_297_itm_17_2_1[15:1])
      + conv_s2s_13_16({Accum2_acc_1586_nl , (input_1_rsci_idat[123:116])}) + conv_s2s_13_16(input_1_rsci_idat[47:35]);
  assign Accum2_acc_768_nl = nl_Accum2_acc_768_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1 = Accum2_acc_769_nl
      + Accum2_acc_768_nl + Accum2_acc_766_cse_1 + Product2_acc_217_itm_17_2_1 +
      Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_777_nl = conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_478_itm_17_2_1[15:2]) + conv_s2s_12_16(input_1_rsci_idat[175:164])
      + conv_s2s_12_16(input_1_rsci_idat[191:180]) + conv_s2s_13_16({Accum2_Accum2_conc_115_12_7
      , (input_1_rsci_idat[202:196])}) + conv_s2s_12_16(input_1_rsci_idat[95:84]);
  assign Accum2_acc_777_nl = nl_Accum2_acc_777_nl[15:0];
  assign nl_Accum2_acc_779_nl = Accum2_acc_777_nl + Product2_acc_152_itm_17_2_1;
  assign Accum2_acc_779_nl = nl_Accum2_acc_779_nl[15:0];
  assign nl_Accum2_acc_778_nl = Product2_acc_238_itm_17_2_1 + Product2_acc_932_itm_19_4_1;
  assign Accum2_acc_778_nl = nl_Accum2_acc_778_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1 = Accum2_acc_779_nl
      + Accum2_acc_778_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1588_nl = conv_s2s_7_8(input_1_rsci_idat[47:41]) + 8'b11111011;
  assign Accum2_acc_1588_nl = nl_Accum2_acc_1588_nl[7:0];
  assign nl_Accum2_acc_787_nl = Accum2_acc_1648 + conv_s2s_15_16(input_1_rsci_idat[223:209])
      + conv_s2s_14_16({Accum2_acc_1588_nl , (input_1_rsci_idat[40:35])}) + conv_s2s_14_16(input_1_rsci_idat[31:18]);
  assign Accum2_acc_787_nl = nl_Accum2_acc_787_nl[15:0];
  assign nl_Accum2_acc_786_nl = Product2_acc_11_itm_17_2_1 + Product2_acc_299_itm_19_4_1;
  assign Accum2_acc_786_nl = nl_Accum2_acc_786_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1 = Accum2_acc_787_nl
      + Accum2_acc_786_nl + Product2_acc_379_itm_18_3_1 + Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_802_itm_17_2_1 + Product2_acc_901_itm_19_4_1;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[14:10]!=5'b00000);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_238_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1
      + conv_s2s_10_13({9'b101100000 , (~ (input_1_rsci_idat[0]))});
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_238_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_238_nl[12:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_246_nl = Product2_acc_871_itm_17_2_1
      + Product2_acc_932_itm_19_4_1 + conv_s2s_15_16(Product2_acc_1086_itm_16_1_1[15:1])
      + conv_s2s_14_16(Product2_acc_122_itm_17_2_1[15:2]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_238_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_246_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_246_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_245_nl = Product2_acc_75_itm_19_4_1
      + conv_s2s_15_16(~ (input_1_rsci_idat[15:1])) + conv_s2s_15_16(Product2_acc_379_itm_18_3_1[15:1]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_245_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_245_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_244_nl = Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_298_itm_17_2_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_244_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_244_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_243_nl = Product2_acc_541_itm_19_4_1
      + Product2_acc_797_cse_sva_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_243_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_243_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_246_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_245_nl + nnet_product_mult_input_t_config2_weight_t_product_acc_244_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_243_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_791_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[63:52]);
  assign Accum2_acc_791_nl = nl_Accum2_acc_791_nl[12:0];
  assign nl_Accum2_acc_1589_nl = conv_s2s_6_7(input_1_rsci_idat[95:90]) + 7'b0000001;
  assign Accum2_acc_1589_nl = nl_Accum2_acc_1589_nl[6:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1 = Product2_acc_601_itm_19_4_1
      + Product2_acc_952_itm_19_4_1 + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_671_itm_18_3_1[15:1]) + conv_s2s_14_16(input_1_rsci_idat[79:66])
      + conv_s2s_14_16(input_1_rsci_idat[111:98]) + conv_s2s_13_16(Accum2_acc_791_nl)
      + conv_s2s_13_16({Accum2_acc_1589_nl , (input_1_rsci_idat[89:84])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[47:35]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_811_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1]);
  assign Accum2_acc_811_nl = nl_Accum2_acc_811_nl[15:0];
  assign nl_Accum2_acc_1590_nl = conv_s2s_4_5(input_1_rsci_idat[207:204]) + 5'b11111;
  assign Accum2_acc_1590_nl = nl_Accum2_acc_1590_nl[4:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1 = Accum2_acc_811_nl
      + conv_s2s_15_16(Accum2_acc_457_cse_1) + conv_s2s_15_16(Product2_acc_1147_itm_16_2_1)
      + conv_s2s_14_16(Product2_acc_532_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2])
      + conv_s2s_13_16({Accum2_acc_1590_nl , (input_1_rsci_idat[203:196])}) + conv_s2s_13_16(input_1_rsci_idat[15:3])
      + conv_s2s_13_16(input_1_rsci_idat[143:131]) + conv_s2s_12_16(input_1_rsci_idat[47:36]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_820_nl = conv_s2s_15_16(Product2_acc_876_itm_18_3_1[15:1])
      + conv_s2s_15_16(input_1_rsci_idat[31:17]) + conv_s2s_15_16(Product2_acc_458_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_216_itm_18_3_1[15:1]);
  assign Accum2_acc_820_nl = nl_Accum2_acc_820_nl[15:0];
  assign nl_Accum2_acc_818_nl = Product2_acc_285_itm_19_4_1 + Product2_acc_1080_itm_16_1_1;
  assign Accum2_acc_818_nl = nl_Accum2_acc_818_nl[15:0];
  assign nl_Accum2_acc_817_nl = Product2_acc_671_itm_18_3_1 + Product2_acc_743_cse_sva_1;
  assign Accum2_acc_817_nl = nl_Accum2_acc_817_nl[15:0];
  assign nl_Accum2_acc_816_nl = Product2_acc_952_itm_19_4_1 + conv_s2s_15_16(Product2_acc_801_itm_18_4_1);
  assign Accum2_acc_816_nl = nl_Accum2_acc_816_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1 = Accum2_acc_820_nl
      + Accum2_acc_818_nl + Product2_acc_154_itm_19_4_1 + Accum2_acc_817_nl + Accum2_acc_816_nl
      + conv_s2s_15_16(Product2_acc_33_itm_15_1_1) + conv_s2s_13_16(input_1_rsci_idat[127:115]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1 = (Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1591_nl = conv_s2s_5_6(input_1_rsci_idat[111:107]) + 6'b111001;
  assign Accum2_acc_1591_nl = nl_Accum2_acc_1591_nl[5:0];
  assign nl_Accum2_acc_833_nl = Product2_acc_951_itm_19_4_1 + conv_s2s_13_16(Accum2_acc_825_cse_1)
      + conv_s2s_13_16({Accum2_acc_1591_nl , (input_1_rsci_idat[106:100])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1);
  assign Accum2_acc_833_nl = nl_Accum2_acc_833_nl[15:0];
  assign nl_Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1 = Accum2_acc_833_nl + conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1])
      + conv_s2s_14_16(input_1_rsci_idat[95:82]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_1064_itm_16_1_1[15:1]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1);
  assign Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1 = (Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_844_nl = conv_s2s_15_16(Product2_acc_796_itm_18_4_1) + conv_s2s_15_16(Product2_acc_604_itm_18_3_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[207:194]) + conv_s2s_14_16(Product2_acc_124_cse_sva_1[15:2]);
  assign Accum2_acc_844_nl = nl_Accum2_acc_844_nl[15:0];
  assign nl_Accum2_acc_843_nl = Product2_acc_1072_itm_17_2_1 + Product2_acc_450_itm_19_4_1;
  assign Accum2_acc_843_nl = nl_Accum2_acc_843_nl[15:0];
  assign nl_Accum2_acc_837_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_123_12_7 , (input_1_rsci_idat[154:148])});
  assign Accum2_acc_837_nl = nl_Accum2_acc_837_nl[13:0];
  assign nl_Accum2_acc_842_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(Accum2_acc_837_nl) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[95:83]);
  assign Accum2_acc_842_nl = nl_Accum2_acc_842_nl[15:0];
  assign nl_Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1 = Accum2_acc_844_nl + Accum2_acc_843_nl
      + Accum2_acc_842_nl;
  assign Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1 = (Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1593_nl = conv_s2s_6_7(input_1_rsci_idat[175:170]) + 7'b1111011;
  assign Accum2_acc_1593_nl = nl_Accum2_acc_1593_nl[6:0];
  assign nl_Accum2_acc_856_nl = conv_s2s_15_16(Product2_acc_796_itm_18_4_1) + conv_s2s_15_16(Product2_acc_538_cse_sva_1[15:1])
      + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_1332_itm_17_2_1[15:2]) + conv_s2s_13_16({Accum2_acc_1593_nl
      , (input_1_rsci_idat[169:164])});
  assign Accum2_acc_856_nl = nl_Accum2_acc_856_nl[15:0];
  assign nl_Accum2_acc_855_nl = Product2_acc_283_itm_18_3_1 + conv_s2s_15_16(Product2_acc_382_cse_sva_1[15:1])
      + conv_s2s_14_16(Accum2_acc_635_cse_1);
  assign Accum2_acc_855_nl = nl_Accum2_acc_855_nl[15:0];
  assign nl_Accum2_acc_854_nl = Product2_acc_476_itm_19_4_1 + conv_s2s_14_16(Product2_acc_871_itm_17_2_1[15:2])
      + conv_s2s_14_16(Product2_acc_943_cse_sva_1[15:2]);
  assign Accum2_acc_854_nl = nl_Accum2_acc_854_nl[15:0];
  assign nl_Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1 = Accum2_acc_856_nl + Accum2_acc_855_nl
      + Accum2_acc_854_nl;
  assign Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1 = (Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1594_nl = conv_s2s_6_7(input_1_rsci_idat[127:122]) + 7'b0000001;
  assign Accum2_acc_1594_nl = nl_Accum2_acc_1594_nl[6:0];
  assign nl_Accum2_acc_863_nl = conv_s2s_15_16(Product2_acc_802_itm_17_2_1[15:1])
      + conv_s2s_14_16(input_1_rsci_idat[143:130]) + conv_s2s_13_16({Accum2_acc_1594_nl
      , (input_1_rsci_idat[121:116])});
  assign Accum2_acc_863_nl = nl_Accum2_acc_863_nl[15:0];
  assign nl_Accum2_acc_867_nl = Accum2_acc_863_nl + Product2_acc_298_itm_17_2_1;
  assign Accum2_acc_867_nl = nl_Accum2_acc_867_nl[15:0];
  assign nl_Accum2_acc_862_nl = (Product2_acc_728_itm_18_3_1[15:1]) + conv_s2s_13_15(input_1_rsci_idat[47:35])
      + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_862_nl = nl_Accum2_acc_862_nl[14:0];
  assign nl_Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1 = Accum2_acc_867_nl + Product2_acc_664_itm_19_4_1
      + Product2_acc_952_itm_19_4_1 + Product2_acc_377_itm_17_2_1 + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Accum2_acc_862_nl) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[63:50]);
  assign Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1 = (Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_876_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(input_1_rsci_idat[207:194]) + conv_s2s_14_16(Product2_acc_629_itm_17_3_1[14:1]);
  assign Accum2_acc_876_nl = nl_Accum2_acc_876_nl[15:0];
  assign nl_Accum2_acc_1595_nl = conv_s2s_6_7(input_1_rsci_idat[63:58]) + 7'b1111111;
  assign Accum2_acc_1595_nl = nl_Accum2_acc_1595_nl[6:0];
  assign nl_Accum2_acc_880_nl = Accum2_acc_876_nl + conv_s2s_15_16(input_1_rsci_idat[47:33])
      + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2]) + conv_s2s_13_16({Accum2_acc_1595_nl
      , (input_1_rsci_idat[57:52])});
  assign Accum2_acc_880_nl = nl_Accum2_acc_880_nl[15:0];
  assign nl_Accum2_acc_879_nl = conv_s2s_15_16(Product2_acc_560_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_283_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_3_itm_15_1_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_879_nl = nl_Accum2_acc_879_nl[15:0];
  assign nl_Accum2_acc_878_nl = Product2_acc_492_itm_17_2_1 + Product2_acc_670_itm_19_4_1;
  assign Accum2_acc_878_nl = nl_Accum2_acc_878_nl[15:0];
  assign nl_Accum2_acc_877_nl = Product2_acc_733_itm_17_2_1 + Product2_acc_795_itm_17_2_1;
  assign Accum2_acc_877_nl = nl_Accum2_acc_877_nl[15:0];
  assign nl_Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1 = Accum2_acc_880_nl + Accum2_acc_879_nl
      + Accum2_acc_878_nl + Accum2_acc_877_nl;
  assign Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1 = (Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_893_nl = Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_379_itm_18_3_1[15:1]) + conv_s2s_14_16(Product2_acc_532_cse_sva_1[15:2])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1);
  assign Accum2_acc_893_nl = nl_Accum2_acc_893_nl[15:0];
  assign nl_Accum2_acc_892_nl = Product2_acc_141_itm_19_4_1 + Product2_acc_298_itm_17_2_1;
  assign Accum2_acc_892_nl = nl_Accum2_acc_892_nl[15:0];
  assign nl_Accum2_acc_1596_nl = conv_s2s_6_7(input_1_rsci_idat[159:154]) + 7'b0000011;
  assign Accum2_acc_1596_nl = nl_Accum2_acc_1596_nl[6:0];
  assign nl_Accum2_acc_890_nl = Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_16({Accum2_acc_1596_nl , (input_1_rsci_idat[153:148])}) + conv_s2s_13_16(input_1_rsci_idat[15:3])
      + conv_s2s_13_16(input_1_rsci_idat[207:195]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1);
  assign Accum2_acc_890_nl = nl_Accum2_acc_890_nl[15:0];
  assign nl_Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1 = Accum2_acc_893_nl + Accum2_acc_892_nl
      + Accum2_acc_890_nl + Product2_acc_478_itm_17_2_1 + Product2_acc_802_itm_17_2_1;
  assign Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1 = (Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_905_nl = conv_s2s_15_16(Product2_acc_1086_itm_16_1_1[15:1])
      + conv_s2s_15_16(Product2_acc_1334_itm_17_3_1) + conv_s2s_15_16(Product2_acc_1336_itm_18_3_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_905_nl = nl_Accum2_acc_905_nl[15:0];
  assign nl_Accum2_acc_1597_nl = conv_s2s_7_8(input_1_rsci_idat[63:57]) + 8'b00000111;
  assign Accum2_acc_1597_nl = nl_Accum2_acc_1597_nl[7:0];
  assign nl_Accum2_acc_898_nl = conv_s2s_15_16(Product2_acc_91_itm_15_1_1) + conv_s2s_14_16({Accum2_acc_1597_nl
      , (input_1_rsci_idat[56:51])});
  assign Accum2_acc_898_nl = nl_Accum2_acc_898_nl[15:0];
  assign nl_Accum2_acc_904_nl = Accum2_acc_898_nl + Product2_acc_1028_itm_17_2_1;
  assign Accum2_acc_904_nl = nl_Accum2_acc_904_nl[15:0];
  assign Product2_acc_1324_nl =  -conv_s2s_12_13(input_1_rsci_idat[47:36]);
  assign nl_Product2_acc_1273_nl = ({(input_1_rsci_idat[47:32]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1324_nl
      , (~ (input_1_rsci_idat[35:32]))});
  assign Product2_acc_1273_nl = nl_Product2_acc_1273_nl[17:0];
  assign nl_Product2_acc_157_nl = conv_s2s_18_20(Product2_acc_1273_nl) + ({(~ (input_1_rsci_idat[47:32]))
      , 4'b0000});
  assign Product2_acc_157_nl = nl_Product2_acc_157_nl[19:0];
  assign nl_Accum2_acc_902_nl = Product2_acc_691_itm_19_4_1 + Product2_acc_794_cse_sva_1;
  assign Accum2_acc_902_nl = nl_Accum2_acc_902_nl[15:0];
  assign nl_Accum2_acc_901_nl = Product2_acc_954_itm_19_4_1 + conv_s2s_14_16(input_1_rsci_idat[207:194])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_901_nl = nl_Accum2_acc_901_nl[15:0];
  assign nl_Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1 = Accum2_acc_905_nl + Accum2_acc_904_nl
      + (readslicef_20_16_4(Product2_acc_157_nl)) + Product2_acc_604_itm_18_3_1 +
      Accum2_acc_902_nl + Accum2_acc_901_nl;
  assign Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1 = (Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_913_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_195_cse_sva_1[15:1]);
  assign Accum2_acc_913_nl = nl_Accum2_acc_913_nl[15:0];
  assign nl_Accum2_acc_916_nl = Accum2_acc_913_nl + Product2_acc_308_cse_sva_1;
  assign Accum2_acc_916_nl = nl_Accum2_acc_916_nl[15:0];
  assign nl_Accum2_acc_910_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_123_12_7 , (input_1_rsci_idat[154:148])});
  assign Accum2_acc_910_nl = nl_Accum2_acc_910_nl[13:0];
  assign nl_Accum2_acc_915_nl = Product2_acc_455_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_910_nl)
      + conv_s2s_14_16(Product2_acc_730_cse_sva_1[15:2]);
  assign Accum2_acc_915_nl = nl_Accum2_acc_915_nl[15:0];
  assign nl_Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1 = Accum2_acc_916_nl + Accum2_acc_915_nl
      + conv_s2s_15_16(Product2_acc_943_cse_sva_1[15:1]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1 = (Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1599_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[12:7])
      + 6'b111101;
  assign Accum2_acc_1599_nl = nl_Accum2_acc_1599_nl[5:0];
  assign nl_Accum2_acc_928_nl = conv_s2s_15_16(Accum2_acc_343_cse_1) + conv_s2s_15_16(Product2_acc_458_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_72_itm_18_3_1[15:1]) + conv_s2s_14_16(Accum2_acc_534_cse_1)
      + conv_s2s_13_16({Accum2_acc_1599_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[6:0])})
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign Accum2_acc_928_nl = nl_Accum2_acc_928_nl[15:0];
  assign nl_Accum2_acc_926_nl = Product2_acc_1079_itm_16_1_1 + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_926_nl = nl_Accum2_acc_926_nl[15:0];
  assign nl_Accum2_acc_925_nl = Product2_acc_1117_itm_16_1_1 + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_925_nl = nl_Accum2_acc_925_nl[15:0];
  assign nl_Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1 = Accum2_acc_928_nl + Accum2_acc_926_nl
      + Accum2_acc_925_nl + Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_330_itm_19_4_1;
  assign Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1 = (Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_933_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_119_12_6 , (input_1_rsci_idat[137:132])});
  assign Accum2_acc_933_nl = nl_Accum2_acc_933_nl[13:0];
  assign nl_Accum2_acc_940_nl = conv_s2s_15_16(Product2_acc_1336_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_1053_itm_16_1_1[15:1]) + conv_s2s_14_16(Accum2_acc_933_nl)
      + conv_s2s_14_16(input_1_rsci_idat[223:210]) + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2]);
  assign Accum2_acc_940_nl = nl_Accum2_acc_940_nl[15:0];
  assign nl_Accum2_acc_935_nl = conv_s2s_14_15(Product2_acc_867_cse_sva_1[15:2])
      + conv_s2s_13_15(input_1_rsci_idat[47:35]) + conv_s2s_13_15(input_1_rsci_idat[127:115]);
  assign Accum2_acc_935_nl = nl_Accum2_acc_935_nl[14:0];
  assign nl_Accum2_acc_938_nl = Product2_acc_742_itm_17_2_1 + conv_s2s_15_16(Accum2_acc_935_nl);
  assign Accum2_acc_938_nl = nl_Accum2_acc_938_nl[15:0];
  assign nl_Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1 = Accum2_acc_940_nl + Accum2_acc_938_nl
      + Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_691_itm_19_4_1;
  assign Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1 = (Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1601_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[12:6])
      + 7'b1110111;
  assign Accum2_acc_1601_nl = nl_Accum2_acc_1601_nl[6:0];
  assign nl_Accum2_acc_944_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1601_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[5:0])});
  assign Accum2_acc_944_nl = nl_Accum2_acc_944_nl[13:0];
  assign nl_Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1 = Accum2_acc_590_cse_1 +
      Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(Accum2_acc_944_nl) + conv_s2s_14_16(input_1_rsci_idat[63:50])
      + conv_s2s_14_16(input_1_rsci_idat[143:130]) + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_934_itm_17_2_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[175:163]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1 = (Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1602_nl = conv_s2s_5_6(input_1_rsci_idat[207:203]) + 6'b111111;
  assign Accum2_acc_1602_nl = nl_Accum2_acc_1602_nl[5:0];
  assign nl_Accum2_acc_958_nl = conv_s2s_14_15(Product2_acc_532_cse_sva_1[15:2])
      + conv_s2s_13_15(Accum2_acc_306_cse_1) + conv_s2s_13_15({Accum2_acc_1602_nl
      , (input_1_rsci_idat[202:196])});
  assign Accum2_acc_958_nl = nl_Accum2_acc_958_nl[14:0];
  assign nl_Accum2_acc_961_nl = Product2_acc_936_cse_sva_1 + conv_s2s_15_16(Accum2_acc_958_nl);
  assign Accum2_acc_961_nl = nl_Accum2_acc_961_nl[15:0];
  assign nl_Accum2_acc_964_nl = Accum2_acc_961_nl + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_308_cse_sva_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_964_nl = nl_Accum2_acc_964_nl[15:0];
  assign nl_Accum2_acc_963_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_665_cse_sva_1[15:1]) + conv_s2s_15_16(Product2_acc_1118_itm_16_1_1[15:1]);
  assign Accum2_acc_963_nl = nl_Accum2_acc_963_nl[15:0];
  assign nl_Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1 = Accum2_acc_964_nl + Accum2_acc_963_nl
      + Product2_acc_367_itm_19_4_1 + Product2_acc_476_itm_19_4_1;
  assign Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1 = (Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_973_nl = Product2_acc_728_itm_18_3_1 + conv_s2s_14_16(Product2_acc_867_cse_sva_1[15:2])
      + conv_s2s_14_16(Product2_acc_532_cse_sva_1[15:2]);
  assign Accum2_acc_973_nl = nl_Accum2_acc_973_nl[15:0];
  assign nl_Accum2_acc_976_nl = Accum2_acc_973_nl + conv_s2s_15_16(Product2_acc_801_itm_18_4_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2]);
  assign Accum2_acc_976_nl = nl_Accum2_acc_976_nl[15:0];
  assign nl_Accum2_acc_975_nl = conv_s2s_15_16(Product2_acc_671_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_970_cse_sva_1[15:1]) + conv_s2s_15_16(Product2_acc_283_itm_18_3_1[15:1])
      + conv_s2s_15_16(input_1_rsci_idat[47:33]);
  assign Accum2_acc_975_nl = nl_Accum2_acc_975_nl[15:0];
  assign nl_Accum2_acc_1603_nl = (Product2_acc_1338_itm_17_3_1[14:7]) + 8'b11111011;
  assign Accum2_acc_1603_nl = nl_Accum2_acc_1603_nl[7:0];
  assign nl_Accum2_acc_974_nl = Product2_acc_476_itm_19_4_1 + conv_s2s_15_16(Product2_acc_1034_itm_16_1_1[15:1])
      + conv_s2s_14_16({Accum2_acc_1603_nl , (Product2_acc_1338_itm_17_3_1[6:1])});
  assign Accum2_acc_974_nl = nl_Accum2_acc_974_nl[15:0];
  assign nl_Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1 = Accum2_acc_976_nl + Accum2_acc_975_nl
      + Accum2_acc_974_nl;
  assign Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1 = (Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_979_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[47:36]);
  assign Accum2_acc_979_nl = nl_Accum2_acc_979_nl[12:0];
  assign nl_Accum2_acc_981_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(Accum2_acc_979_nl);
  assign Accum2_acc_981_nl = nl_Accum2_acc_981_nl[13:0];
  assign nl_Accum2_acc_988_nl = conv_s2s_15_16(Product2_acc_728_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_499_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_379_itm_18_3_1[15:1])
      + conv_s2s_14_16(Accum2_acc_981_nl);
  assign Accum2_acc_988_nl = nl_Accum2_acc_988_nl[15:0];
  assign nl_Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1 = Accum2_acc_988_nl + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_691_itm_19_4_1 + Product2_acc_216_itm_18_3_1 + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_867_cse_sva_1[15:1]) + conv_s2s_14_16(Product2_acc_3_itm_15_1_1[14:1])
      + conv_s2s_13_16({Accum2_Accum2_conc_121_12_8 , (input_1_rsci_idat[219:212])})
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1);
  assign Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1 = (Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1000_nl = Product2_acc_601_itm_19_4_1 + conv_s2s_15_16(Product2_acc_1086_itm_16_1_1[15:1])
      + conv_s2s_14_16(Product2_acc_217_itm_17_2_1[15:2]) + conv_s2s_13_16(Accum2_acc_532_cse_1);
  assign Accum2_acc_1000_nl = nl_Accum2_acc_1000_nl[15:0];
  assign nl_Accum2_acc_995_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15(Accum2_acc_992_cse_1);
  assign Accum2_acc_995_nl = nl_Accum2_acc_995_nl[14:0];
  assign nl_Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1000_nl + Product2_acc_834_itm_19_4_1
      + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_769_itm_19_4_1 + conv_s2s_15_16(Accum2_acc_995_nl) + conv_s2s_14_16(Product2_acc_934_itm_17_2_1[15:2])
      + conv_s2s_14_16(input_1_rsci_idat[79:66]);
  assign Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1 = (Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1013_nl = conv_s2s_15_16(Product2_acc_946_itm_18_3_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_1042_itm_16_1_1[15:1]) + conv_s2s_15_16(Product2_acc_62_itm_18_4_1);
  assign Accum2_acc_1013_nl = nl_Accum2_acc_1013_nl[15:0];
  assign Product2_acc_1325_nl =  -conv_s2s_13_14(input_1_rsci_idat[143:131]);
  assign nl_Product2_acc_644_nl = conv_s2s_17_20({Product2_acc_1325_nl , (~ (input_1_rsci_idat[130:128]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[143:128])) , 3'b001});
  assign Product2_acc_644_nl = nl_Product2_acc_644_nl[19:0];
  assign nl_Accum2_acc_1012_nl = (readslicef_20_16_4(Product2_acc_644_nl)) + conv_s2s_14_16(input_1_rsci_idat[111:98])
      + conv_s2s_13_16({Accum2_Accum2_conc_117_12_6 , (input_1_rsci_idat[201:196])})
      + conv_s2s_12_16(input_1_rsci_idat[63:52]);
  assign Accum2_acc_1012_nl = nl_Accum2_acc_1012_nl[15:0];
  assign nl_Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1013_nl + Accum2_acc_1012_nl
      + conv_s2s_14_16(input_1_rsci_idat[175:162]) + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2])
      + conv_s2s_14_16(Product2_acc_1338_itm_17_3_1[14:1]) + conv_s2s_12_16(input_1_rsci_idat[79:68])
      + conv_s2s_12_16(input_1_rsci_idat[159:148]);
  assign Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1 = (Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1606_nl = conv_s2s_7_8(input_1_rsci_idat[175:169]) + 8'b00000011;
  assign Accum2_acc_1606_nl = nl_Accum2_acc_1606_nl[7:0];
  assign nl_Accum2_acc_1023_nl = conv_s2s_15_16(Product2_acc_1147_itm_16_2_1) + conv_s2s_13_16(input_1_rsci_idat[15:3])
      + conv_s2s_13_16(input_1_rsci_idat[79:67]) + conv_s2s_14_16({Accum2_acc_1606_nl
      , (input_1_rsci_idat[168:163])}) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[31:18]) + conv_s2s_14_16(input_1_rsci_idat[111:98]);
  assign Accum2_acc_1023_nl = nl_Accum2_acc_1023_nl[15:0];
  assign nl_Accum2_acc_1022_nl = Product2_acc_154_itm_19_4_1 + Product2_acc_547_itm_17_2_1;
  assign Accum2_acc_1022_nl = nl_Accum2_acc_1022_nl[15:0];
  assign nl_Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1023_nl + Accum2_acc_1022_nl
      + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_901_itm_19_4_1;
  assign Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1 = (Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1033_nl = Product2_acc_492_itm_17_2_1 + Product2_acc_942_itm_17_2_1;
  assign Accum2_acc_1033_nl = nl_Accum2_acc_1033_nl[15:0];
  assign nl_Accum2_acc_1032_nl = conv_s2s_14_16(Accum2_acc_1028_cse_1) + conv_s2s_14_16(Accum2_acc_1027_cse_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[127:115]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_1032_nl = nl_Accum2_acc_1032_nl[15:0];
  assign nl_Accum2_acc_1035_nl = Accum2_acc_1033_nl + Accum2_acc_1032_nl;
  assign Accum2_acc_1035_nl = nl_Accum2_acc_1035_nl[15:0];
  assign nl_Accum2_acc_1031_nl = conv_s2s_15_16(Product2_acc_871_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_217_itm_17_2_1[15:1]);
  assign Accum2_acc_1031_nl = nl_Accum2_acc_1031_nl[15:0];
  assign nl_Accum2_acc_1034_nl = Accum2_acc_1031_nl + Product2_acc_1079_itm_16_1_1;
  assign Accum2_acc_1034_nl = nl_Accum2_acc_1034_nl[15:0];
  assign nl_Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1035_nl + Accum2_acc_1034_nl;
  assign Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1 = (Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1046_nl = Product2_acc_1064_itm_16_1_1 + Product2_acc_970_cse_sva_1;
  assign Accum2_acc_1046_nl = nl_Accum2_acc_1046_nl[15:0];
  assign nl_Accum2_acc_1038_nl = (Product2_acc_1332_itm_17_2_1[15:2]) + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign Accum2_acc_1038_nl = nl_Accum2_acc_1038_nl[13:0];
  assign nl_Accum2_acc_1608_nl = conv_s2s_6_7(input_1_rsci_idat[95:90]) + 7'b1111011;
  assign Accum2_acc_1608_nl = nl_Accum2_acc_1608_nl[6:0];
  assign nl_Accum2_acc_1045_nl = conv_s2s_14_16(Accum2_acc_1038_nl) + conv_s2s_14_16({Accum2_acc_1608_nl
      , (input_1_rsci_idat[89:83])}) + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1);
  assign Accum2_acc_1045_nl = nl_Accum2_acc_1045_nl[15:0];
  assign nl_Accum2_acc_1048_nl = Accum2_acc_1046_nl + Accum2_acc_1045_nl;
  assign Accum2_acc_1048_nl = nl_Accum2_acc_1048_nl[15:0];
  assign nl_Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1048_nl + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_532_cse_sva_1[15:2]) + conv_s2s_15_16(Product2_acc_478_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_195_cse_sva_1[15:1]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1 = (Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1058_nl = Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_887_itm_15_1_1) + conv_s2s_15_16(Product2_acc_1334_itm_17_3_1);
  assign Accum2_acc_1058_nl = nl_Accum2_acc_1058_nl[15:0];
  assign nl_Accum2_acc_1609_nl = conv_s2s_6_7(input_1_rsci_idat[143:138]) + 7'b0001001;
  assign Accum2_acc_1609_nl = nl_Accum2_acc_1609_nl[6:0];
  assign nl_Accum2_acc_1054_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_15({Accum2_acc_1609_nl , (input_1_rsci_idat[137:132])}) + conv_s2s_12_15(input_1_rsci_idat[31:20])
      + conv_s2s_12_15(input_1_rsci_idat[47:36]);
  assign Accum2_acc_1054_nl = nl_Accum2_acc_1054_nl[14:0];
  assign nl_Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1058_nl + Product2_acc_455_itm_19_4_1
      + Product2_acc_954_itm_19_4_1 + conv_s2s_15_16(Accum2_acc_1054_nl) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[95:83]);
  assign Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1 = (Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1610_nl = conv_s2s_5_6(input_1_rsci_idat[15:11]) + 6'b111111;
  assign Accum2_acc_1610_nl = nl_Accum2_acc_1610_nl[5:0];
  assign nl_Accum2_acc_1064_nl = conv_s2s_14_15(input_1_rsci_idat[127:114]) + conv_s2s_13_15({Accum2_acc_1610_nl
      , (input_1_rsci_idat[10:4])}) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1);
  assign Accum2_acc_1064_nl = nl_Accum2_acc_1064_nl[14:0];
  assign nl_Accum2_acc_1068_nl = Product2_acc_1144_itm_16_1_1 + conv_s2s_15_16(Accum2_acc_1064_nl);
  assign Accum2_acc_1068_nl = nl_Accum2_acc_1068_nl[15:0];
  assign nl_Accum2_acc_1071_nl = Accum2_acc_1068_nl + conv_s2s_14_16(input_1_rsci_idat[207:194])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_122_itm_17_2_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1071_nl = nl_Accum2_acc_1071_nl[15:0];
  assign nl_Accum2_acc_1070_nl = Accum2_acc_1066_cse_1 + conv_s2s_15_16(Product2_acc_792_cse_sva_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1070_nl = nl_Accum2_acc_1070_nl[15:0];
  assign nl_Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1071_nl + Accum2_acc_1070_nl
      + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_727_itm_19_4_1;
  assign Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1 = (Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign Product2_acc_1326_nl =  -conv_s2s_12_13(input_1_rsci_idat[15:4]);
  assign nl_Product2_acc_1276_nl = ({(input_1_rsci_idat[15:0]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1326_nl
      , (~ (input_1_rsci_idat[3:0]))});
  assign Product2_acc_1276_nl = nl_Product2_acc_1276_nl[17:0];
  assign nl_Product2_acc_41_nl = conv_s2s_18_20(Product2_acc_1276_nl) + ({(~ (input_1_rsci_idat[15:0]))
      , 4'b0000});
  assign Product2_acc_41_nl = nl_Product2_acc_41_nl[19:0];
  assign nl_Accum2_acc_1081_nl = (readslicef_20_16_4(Product2_acc_41_nl)) + Product2_acc_1042_itm_16_1_1;
  assign Accum2_acc_1081_nl = nl_Accum2_acc_1081_nl[15:0];
  assign nl_Accum2_acc_1080_nl = Product2_acc_191_itm_19_4_1 + Product2_acc_394_itm_17_2_1;
  assign Accum2_acc_1080_nl = nl_Accum2_acc_1080_nl[15:0];
  assign nl_Accum2_acc_1084_nl = Accum2_acc_1081_nl + Accum2_acc_1080_nl;
  assign Accum2_acc_1084_nl = nl_Accum2_acc_1084_nl[15:0];
  assign nl_Accum2_acc_1082_nl = conv_s2s_15_16(Product2_acc_943_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_1110_itm_16_2_1) + conv_s2s_15_16(Product2_acc_538_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_297_itm_17_2_1[15:1]);
  assign Accum2_acc_1082_nl = nl_Accum2_acc_1082_nl[15:0];
  assign nl_Accum2_acc_1611_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1[12:6])
      + 7'b1111111;
  assign Accum2_acc_1611_nl = nl_Accum2_acc_1611_nl[6:0];
  assign nl_Accum2_acc_1075_nl = conv_s2s_14_15(Product2_acc_85_itm_15_1_1[14:1])
      + conv_s2s_13_15({Accum2_acc_1611_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1[5:0])})
      + conv_s2s_13_15(input_1_rsci_idat[207:195]);
  assign Accum2_acc_1075_nl = nl_Accum2_acc_1075_nl[14:0];
  assign nl_Accum2_acc_1078_nl = Product2_acc_1125_itm_16_1_1 + conv_s2s_15_16(Accum2_acc_1075_nl);
  assign Accum2_acc_1078_nl = nl_Accum2_acc_1078_nl[15:0];
  assign nl_Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1084_nl + Accum2_acc_1082_nl
      + Accum2_acc_1078_nl + Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_772_itm_18_3_1;
  assign Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1 = (Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1612_nl = conv_s2s_6_7(Product2_acc_370_cse_sva_1[15:10])
      + 7'b0000001;
  assign Accum2_acc_1612_nl = nl_Accum2_acc_1612_nl[6:0];
  assign nl_Accum2_acc_1095_nl = conv_s2s_15_16({Accum2_acc_1612_nl , (Product2_acc_370_cse_sva_1[9:2])})
      + conv_s2s_15_16(Product2_acc_772_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_604_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_1330_itm_17_3_1);
  assign Accum2_acc_1095_nl = nl_Accum2_acc_1095_nl[15:0];
  assign nl_Accum2_acc_1094_nl = conv_s2s_15_16(Product2_acc_308_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_91_itm_15_1_1)
      + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2]);
  assign Accum2_acc_1094_nl = nl_Accum2_acc_1094_nl[15:0];
  assign nl_Accum2_acc_1093_nl = Product2_acc_214_cse_sva_1 + Product2_acc_455_itm_19_4_1;
  assign Accum2_acc_1093_nl = nl_Accum2_acc_1093_nl[15:0];
  assign nl_Accum2_acc_1092_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(input_1_rsci_idat[47:34]) + conv_s2s_14_16(input_1_rsci_idat[127:114]);
  assign Accum2_acc_1092_nl = nl_Accum2_acc_1092_nl[15:0];
  assign nl_Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1095_nl + Accum2_acc_1094_nl
      + Accum2_acc_1093_nl + Accum2_acc_1092_nl;
  assign Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1 = (Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1613_nl = conv_s2s_6_7(input_1_rsci_idat[159:154]) + 7'b1111011;
  assign Accum2_acc_1613_nl = nl_Accum2_acc_1613_nl[6:0];
  assign nl_Accum2_acc_1107_nl = Product2_acc_934_itm_17_2_1 + conv_s2s_13_16({Accum2_acc_1613_nl
      , (input_1_rsci_idat[153:148])}) + conv_s2s_13_16(input_1_rsci_idat[95:83])
      + conv_s2s_13_16(input_1_rsci_idat[111:99]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign Accum2_acc_1107_nl = nl_Accum2_acc_1107_nl[15:0];
  assign nl_Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1107_nl + Product2_acc_1332_itm_17_2_1
      + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2]) + conv_s2s_14_16(Product2_acc_217_itm_17_2_1[15:2])
      + conv_s2s_12_16(input_1_rsci_idat[15:4]) + conv_s2s_12_16(input_1_rsci_idat[79:68])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1);
  assign Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1 = (Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1 = conv_s2s_15_16(Accum2_acc_447_cse_1)
      + conv_s2s_14_16(input_1_rsci_idat[223:210]) + conv_s2s_14_16(Product2_acc_730_cse_sva_1[15:2])
      + conv_s2s_14_16(Product2_acc_802_itm_17_2_1[15:2]) + conv_s2s_14_16(Product2_acc_667_cse_sva_1[15:2])
      + conv_s2s_14_16(Product2_acc_1334_itm_17_3_1[14:1]) + conv_s2s_12_16(input_1_rsci_idat[15:4])
      + conv_s2s_12_16(input_1_rsci_idat[111:100]) + conv_s2s_15_16(Product2_acc_609_cse_sva_1[15:1])
      + conv_s2s_13_16(input_1_rsci_idat[207:195]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1 = (Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1614_nl = conv_s2s_6_7(input_1_rsci_idat[111:106]) + 7'b1111101;
  assign Accum2_acc_1614_nl = nl_Accum2_acc_1614_nl[6:0];
  assign nl_Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1 = Product2_acc_166_itm_18_3_1
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_970_cse_sva_1[15:1]) + conv_s2s_14_16(Product2_acc_297_itm_17_2_1[15:2])
      + conv_s2s_13_16(Accum2_acc_1120_cse_1) + conv_s2s_14_16(input_1_rsci_idat[15:2])
      + conv_s2s_14_16(input_1_rsci_idat[127:114]) + conv_s2s_13_16({Accum2_acc_1614_nl
      , (input_1_rsci_idat[105:100])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1);
  assign Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1 = (Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1138_nl = conv_s2s_15_16(Product2_acc_1147_itm_16_2_1) + conv_s2s_15_16(Product2_acc_217_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_1027_itm_16_2_1) + conv_s2s_14_16(Product2_acc_532_cse_sva_1[15:2])
      + conv_s2s_14_16(Product2_acc_308_cse_sva_1[15:2]);
  assign Accum2_acc_1138_nl = nl_Accum2_acc_1138_nl[15:0];
  assign nl_Accum2_acc_1129_nl = (Product2_acc_122_itm_17_2_1[15:2]) + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1);
  assign Accum2_acc_1129_nl = nl_Accum2_acc_1129_nl[13:0];
  assign nl_Accum2_acc_1137_nl = Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_1034_itm_16_1_1[15:1]) + conv_s2s_14_16(Accum2_acc_1129_nl);
  assign Accum2_acc_1137_nl = nl_Accum2_acc_1137_nl[15:0];
  assign nl_Accum2_acc_1136_nl = Product2_acc_455_itm_19_4_1 + Product2_acc_1105_itm_16_1_1;
  assign Accum2_acc_1136_nl = nl_Accum2_acc_1136_nl[15:0];
  assign nl_Accum2_acc_1615_nl = conv_s2s_7_8(input_1_rsci_idat[159:153]) + 8'b11111101;
  assign Accum2_acc_1615_nl = nl_Accum2_acc_1615_nl[7:0];
  assign nl_Accum2_acc_1131_nl = conv_s2s_14_15({Accum2_acc_1615_nl , (input_1_rsci_idat[152:147])})
      + conv_s2s_14_15(Product2_acc_867_cse_sva_1[15:2]);
  assign Accum2_acc_1131_nl = nl_Accum2_acc_1131_nl[14:0];
  assign nl_Accum2_acc_1135_nl = Product2_acc_1117_itm_16_1_1 + conv_s2s_15_16(Accum2_acc_1131_nl);
  assign Accum2_acc_1135_nl = nl_Accum2_acc_1135_nl[15:0];
  assign nl_Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1138_nl + Accum2_acc_1137_nl
      + Accum2_acc_1136_nl + Accum2_acc_1135_nl;
  assign Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1 = (Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1616_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1[12:6])
      + 7'b0000001;
  assign Accum2_acc_1616_nl = nl_Accum2_acc_1616_nl[6:0];
  assign nl_Accum2_acc_1148_nl = Product2_acc_952_itm_19_4_1 + conv_s2s_15_16(Product2_acc_1042_itm_16_1_1[15:1])
      + conv_s2s_13_16({Accum2_acc_1616_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1[5:0])})
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1);
  assign Accum2_acc_1148_nl = nl_Accum2_acc_1148_nl[15:0];
  assign nl_Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1148_nl + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_297_itm_17_2_1[15:2]) + conv_s2s_15_16(Product2_acc_802_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_1095_itm_16_1_1[15:1]) + conv_s2s_14_16(Product2_acc_377_itm_17_2_1[15:2])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1 = (Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1153_nl = (Product2_acc_934_itm_17_2_1[15:1]) + conv_s2s_14_15(Accum2_acc_295_cse_1);
  assign Accum2_acc_1153_nl = nl_Accum2_acc_1153_nl[14:0];
  assign nl_Accum2_acc_1155_nl = Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Accum2_acc_1153_nl);
  assign Accum2_acc_1155_nl = nl_Accum2_acc_1155_nl[15:0];
  assign nl_Accum2_acc_1617_nl = conv_s2s_6_7(input_1_rsci_idat[143:138]) + 7'b1111001;
  assign Accum2_acc_1617_nl = nl_Accum2_acc_1617_nl[6:0];
  assign nl_Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1155_nl + Product2_acc_281_itm_19_4_1
      + Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_1334_itm_17_3_1) + conv_s2s_14_16(Product2_acc_217_itm_17_2_1[15:2])
      + conv_s2s_13_16({Accum2_acc_1617_nl , (input_1_rsci_idat[137:132])});
  assign Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1 = (Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1159_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[79:68]);
  assign Accum2_acc_1159_nl = nl_Accum2_acc_1159_nl[12:0];
  assign nl_Accum2_acc_1618_nl = conv_s2s_6_7(input_1_rsci_idat[207:202]) + 7'b0000111;
  assign Accum2_acc_1618_nl = nl_Accum2_acc_1618_nl[6:0];
  assign nl_Accum2_acc_1167_nl = conv_s2s_15_16(input_1_rsci_idat[111:97]) + conv_s2s_15_16(Product2_acc_730_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_1332_itm_17_2_1[15:1]) + conv_s2s_13_16(Accum2_acc_1159_nl)
      + conv_s2s_13_16({Accum2_acc_1618_nl , (input_1_rsci_idat[201:196])});
  assign Accum2_acc_1167_nl = nl_Accum2_acc_1167_nl[15:0];
  assign nl_Accum2_acc_1166_nl = Product2_acc_1042_itm_16_1_1 + Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1166_nl = nl_Accum2_acc_1166_nl[15:0];
  assign nl_Accum2_acc_1164_nl = Product2_acc_946_itm_18_3_1 + conv_s2s_14_16(input_1_rsci_idat[191:178])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1164_nl = nl_Accum2_acc_1164_nl[15:0];
  assign nl_Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1167_nl + Accum2_acc_1166_nl
      + Accum2_acc_766_cse_1 + Accum2_acc_1164_nl;
  assign Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1 = (Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1619_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1[12:6])
      + 7'b0001001;
  assign Accum2_acc_1619_nl = nl_Accum2_acc_1619_nl[6:0];
  assign nl_Accum2_acc_1173_nl = Product2_acc_954_itm_19_4_1 + conv_s2s_14_16(Product2_acc_3_itm_15_1_1[14:1])
      + conv_s2s_13_16({Accum2_acc_1619_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1[5:0])});
  assign Accum2_acc_1173_nl = nl_Accum2_acc_1173_nl[15:0];
  assign nl_Accum2_acc_1178_nl = Accum2_acc_1173_nl + conv_s2s_15_16(Product2_acc_1126_itm_16_1_1[15:1])
      + conv_s2s_14_16(input_1_rsci_idat[127:114]);
  assign Accum2_acc_1178_nl = nl_Accum2_acc_1178_nl[15:0];
  assign nl_Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1178_nl + Product2_acc_72_itm_18_3_1
      + Product2_acc_141_itm_19_4_1 + Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_727_itm_19_4_1 + Product2_acc_876_itm_18_3_1 + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_499_itm_18_3_1;
  assign Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1 = (Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1184_nl = (Product2_acc_217_itm_17_2_1[15:2]) + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1);
  assign Accum2_acc_1184_nl = nl_Accum2_acc_1184_nl[13:0];
  assign nl_Accum2_acc_1192_nl = conv_s2s_15_16(Product2_acc_943_cse_sva_1[15:1])
      + conv_s2s_15_16(input_1_rsci_idat[111:97]) + conv_s2s_15_16(Product2_acc_itm_18_3_1[15:1])
      + conv_s2s_14_16(Accum2_acc_1184_nl);
  assign Accum2_acc_1192_nl = nl_Accum2_acc_1192_nl[15:0];
  assign nl_Accum2_acc_1620_nl = conv_s2s_6_7(input_1_rsci_idat[127:122]) + 7'b1111101;
  assign Accum2_acc_1620_nl = nl_Accum2_acc_1620_nl[6:0];
  assign nl_Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1192_nl + conv_s2s_14_16(Accum2_acc_992_cse_1)
      + conv_s2s_14_16({Accum2_acc_1620_nl , (input_1_rsci_idat[121:115])}) + conv_s2s_15_16(Product2_acc_1105_itm_16_1_1[15:1])
      + conv_s2s_14_16(Product2_acc_308_cse_sva_1[15:2]) + conv_s2s_14_16(Product2_acc_122_itm_17_2_1[15:2])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_667_cse_sva_1[15:2]);
  assign Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1 = (Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1199_nl = Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_16({Accum2_Accum2_conc_117_12_6 , (input_1_rsci_idat[201:196])})
      + conv_s2s_13_16(input_1_rsci_idat[79:67]) + conv_s2s_13_16(input_1_rsci_idat[111:99])
      + conv_s2s_13_16(input_1_rsci_idat[175:163]);
  assign Accum2_acc_1199_nl = nl_Accum2_acc_1199_nl[15:0];
  assign nl_Accum2_acc_1203_nl = Accum2_acc_1199_nl + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_665_cse_sva_1[15:1]);
  assign Accum2_acc_1203_nl = nl_Accum2_acc_1203_nl[15:0];
  assign nl_Product2_acc_1277_nl = (~ (input_1_rsci_idat[47:32])) + conv_s2s_14_16(input_1_rsci_idat[47:34]);
  assign Product2_acc_1277_nl = nl_Product2_acc_1277_nl[15:0];
  assign nl_Product2_acc_1050_nl = conv_s2u_16_18(Product2_acc_1277_nl) + ({(input_1_rsci_idat[47:32])
      , 2'b01});
  assign Product2_acc_1050_nl = nl_Product2_acc_1050_nl[17:0];
  assign nl_Accum2_acc_1201_nl = (readslicef_18_16_2(Product2_acc_1050_nl)) + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1201_nl = nl_Accum2_acc_1201_nl[15:0];
  assign nl_Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1203_nl + Accum2_acc_1201_nl
      + Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_528_itm_19_4_1 + Product2_acc_8_itm_18_3_1 + Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1 = (Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1215_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_458_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_212_itm_18_3_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1215_nl = nl_Accum2_acc_1215_nl[15:0];
  assign nl_Accum2_acc_1622_nl = conv_s2s_5_6(input_1_rsci_idat[143:139]) + 6'b111101;
  assign Accum2_acc_1622_nl = nl_Accum2_acc_1622_nl[5:0];
  assign nl_Accum2_acc_1214_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_127_cse_sva_1[15:1]) + conv_s2s_13_16({Accum2_acc_1622_nl
      , (input_1_rsci_idat[138:132])}) + conv_s2s_12_16(input_1_rsci_idat[15:4]);
  assign Accum2_acc_1214_nl = nl_Accum2_acc_1214_nl[15:0];
  assign nl_Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1215_nl + Accum2_acc_1214_nl
      + conv_s2s_14_16(Product2_acc_867_cse_sva_1[15:2]) + conv_s2s_14_16(input_1_rsci_idat[223:210])
      + conv_s2s_14_16(Product2_acc_733_itm_17_2_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1 = (Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1623_nl = conv_s2s_5_6(input_1_rsci_idat[207:203]) + 6'b111101;
  assign Accum2_acc_1623_nl = nl_Accum2_acc_1623_nl[5:0];
  assign nl_Accum2_acc_1220_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1623_nl , (input_1_rsci_idat[202:196])});
  assign Accum2_acc_1220_nl = nl_Accum2_acc_1220_nl[13:0];
  assign nl_Accum2_acc_1225_nl = Product2_acc_531_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_1220_nl)
      + conv_s2s_13_16(input_1_rsci_idat[47:35]) + conv_s2s_13_16(input_1_rsci_idat[175:163]);
  assign Accum2_acc_1225_nl = nl_Accum2_acc_1225_nl[15:0];
  assign nl_Accum2_acc_1228_nl = Accum2_acc_1225_nl + conv_s2s_15_16(Product2_acc_937_itm_18_3_1[15:1])
      + conv_s2s_14_16(Accum2_acc_727_cse_1) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1228_nl = nl_Accum2_acc_1228_nl[15:0];
  assign nl_Accum2_acc_1227_nl = Product2_acc_212_itm_18_3_1 + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_429_itm_18_3_1[15:1]);
  assign Accum2_acc_1227_nl = nl_Accum2_acc_1227_nl[15:0];
  assign nl_Accum2_acc_1226_nl = Product2_acc_1066_itm_16_1_1 + Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1226_nl = nl_Accum2_acc_1226_nl[15:0];
  assign nl_Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1228_nl + Accum2_acc_1227_nl
      + Accum2_acc_1226_nl;
  assign Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1 = (Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign Product2_acc_1327_nl =  -conv_s2s_13_14(input_1_rsci_idat[47:35]);
  assign nl_Product2_acc_174_nl = conv_s2s_17_20({Product2_acc_1327_nl , (~ (input_1_rsci_idat[34:32]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[47:32])) , 3'b001});
  assign Product2_acc_174_nl = nl_Product2_acc_174_nl[19:0];
  assign nl_Accum2_acc_1237_nl = (readslicef_20_16_4(Product2_acc_174_nl)) + Product2_acc_214_cse_sva_1;
  assign Accum2_acc_1237_nl = nl_Accum2_acc_1237_nl[15:0];
  assign nl_Accum2_acc_1236_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1236_nl = nl_Accum2_acc_1236_nl[15:0];
  assign nl_Accum2_acc_1240_nl = Accum2_acc_1237_nl + Accum2_acc_1236_nl;
  assign Accum2_acc_1240_nl = nl_Accum2_acc_1240_nl[15:0];
  assign nl_Accum2_acc_1624_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[12:7])
      + 6'b111111;
  assign Accum2_acc_1624_nl = nl_Accum2_acc_1624_nl[5:0];
  assign nl_Accum2_acc_1238_nl = conv_s2s_15_16(input_1_rsci_idat[31:17]) + conv_s2s_15_16(Product2_acc_728_itm_18_3_1[15:1])
      + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2]) + conv_s2s_14_16(input_1_rsci_idat[207:194])
      + conv_s2s_13_16({Accum2_acc_1624_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[6:0])});
  assign Accum2_acc_1238_nl = nl_Accum2_acc_1238_nl[15:0];
  assign nl_Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1240_nl + Accum2_acc_1238_nl
      + Accum2_acc_426_cse_1 + Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_932_itm_19_4_1;
  assign Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1 = (Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1252_nl = Product2_acc_127_cse_sva_1 + Product2_acc_1072_itm_17_2_1;
  assign Accum2_acc_1252_nl = nl_Accum2_acc_1252_nl[15:0];
  assign nl_Accum2_acc_1251_nl = Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_1086_itm_16_1_1;
  assign Accum2_acc_1251_nl = nl_Accum2_acc_1251_nl[15:0];
  assign nl_Accum2_acc_1254_nl = Accum2_acc_1252_nl + Accum2_acc_1251_nl;
  assign Accum2_acc_1254_nl = nl_Accum2_acc_1254_nl[15:0];
  assign nl_Accum2_acc_1243_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[31:20]);
  assign Accum2_acc_1243_nl = nl_Accum2_acc_1243_nl[12:0];
  assign nl_Accum2_acc_1625_nl = conv_s2s_5_6(input_1_rsci_idat[175:171]) + 6'b111111;
  assign Accum2_acc_1625_nl = nl_Accum2_acc_1625_nl[5:0];
  assign nl_Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1254_nl + conv_s2s_15_16(Product2_acc_797_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_604_itm_18_3_1[15:1]) + conv_s2s_14_16(input_1_rsci_idat[63:50])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1)
      + conv_s2s_13_16(Accum2_acc_1243_nl) + conv_s2s_13_16({Accum2_acc_1625_nl ,
      (input_1_rsci_idat[170:164])}) + conv_s2s_13_16(input_1_rsci_idat[207:195])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1);
  assign Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1 = (Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1264_nl = conv_s2s_15_16(Product2_acc_1147_itm_16_2_1) + conv_s2s_15_16(Product2_acc_671_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_609_cse_sva_1[15:1]) + conv_s2s_15_16(Product2_acc_217_itm_17_2_1[15:1]);
  assign Accum2_acc_1264_nl = nl_Accum2_acc_1264_nl[15:0];
  assign nl_Accum2_acc_1258_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(Accum2_acc_825_cse_1);
  assign Accum2_acc_1258_nl = nl_Accum2_acc_1258_nl[13:0];
  assign nl_Accum2_acc_1262_nl = Product2_acc_809_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_1258_nl)
      + conv_s2s_13_16({Accum2_Accum2_conc_127_12_7 , (input_1_rsci_idat[170:164])})
      + conv_s2s_13_16(input_1_rsci_idat[127:115]);
  assign Accum2_acc_1262_nl = nl_Accum2_acc_1262_nl[15:0];
  assign nl_Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1264_nl + Accum2_acc_1262_nl
      + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_456_itm_19_4_1;
  assign Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1 = (Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1270_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_115_12_7 , (input_1_rsci_idat[202:196])});
  assign Accum2_acc_1270_nl = nl_Accum2_acc_1270_nl[13:0];
  assign nl_Accum2_acc_1276_nl = Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_283_itm_18_3_1[15:1]) + conv_s2s_14_16(Accum2_acc_1270_nl);
  assign Accum2_acc_1276_nl = nl_Accum2_acc_1276_nl[15:0];
  assign nl_Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1276_nl + Accum2_acc_1648
      + conv_s2s_14_16(Accum2_acc_1027_cse_1) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[47:35]) + conv_s2s_13_16(input_1_rsci_idat[223:211]);
  assign Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1 = (Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1628_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[12:6])
      + 7'b1111001;
  assign Accum2_acc_1628_nl = nl_Accum2_acc_1628_nl[6:0];
  assign nl_Accum2_acc_1288_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1]) + conv_s2s_13_16({Accum2_acc_1628_nl
      , (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[5:0])})
      + conv_s2s_13_16(input_1_rsci_idat[31:19]) + conv_s2s_13_16(input_1_rsci_idat[111:99])
      + conv_s2s_13_16(input_1_rsci_idat[143:131]);
  assign Accum2_acc_1288_nl = nl_Accum2_acc_1288_nl[15:0];
  assign nl_Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1288_nl + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[159:146]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_124_cse_sva_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[175:162]) + conv_s2s_14_16(input_1_rsci_idat[207:194]);
  assign Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1 = (Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1297_nl = conv_s2s_15_16(Product2_acc_772_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_802_itm_17_2_1[15:1]) + conv_s2s_15_16(Product2_acc_379_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_458_itm_18_3_1[15:1]);
  assign Accum2_acc_1297_nl = nl_Accum2_acc_1297_nl[15:0];
  assign nl_Accum2_acc_1296_nl = Product2_acc_166_itm_18_3_1 + conv_s2s_15_16(Product2_acc_195_cse_sva_1[15:1])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1296_nl = nl_Accum2_acc_1296_nl[15:0];
  assign nl_Accum2_acc_1629_nl = conv_s2s_8_9(Product2_acc_85_itm_15_1_1[14:7]) +
      9'b000000001;
  assign Accum2_acc_1629_nl = nl_Accum2_acc_1629_nl[8:0];
  assign nl_Accum2_acc_1294_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16({Accum2_acc_1629_nl , (Product2_acc_85_itm_15_1_1[6:1])});
  assign Accum2_acc_1294_nl = nl_Accum2_acc_1294_nl[15:0];
  assign nl_Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1297_nl + Accum2_acc_1296_nl
      + Accum2_acc_1294_nl + Product2_acc_330_itm_19_4_1 + Product2_acc_541_itm_19_4_1;
  assign Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1 = (Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1303_nl = conv_s2s_15_16(Product2_acc_867_cse_sva_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1303_nl = nl_Accum2_acc_1303_nl[15:0];
  assign nl_Accum2_acc_1308_nl = Accum2_acc_1303_nl + Product2_acc_1028_itm_17_2_1;
  assign Accum2_acc_1308_nl = nl_Accum2_acc_1308_nl[15:0];
  assign nl_Accum2_acc_1305_nl = Product2_acc_666_itm_18_3_1 + Product2_acc_1117_itm_16_1_1;
  assign Accum2_acc_1305_nl = nl_Accum2_acc_1305_nl[15:0];
  assign nl_Accum2_acc_1630_nl = conv_s2s_5_6(input_1_rsci_idat[63:59]) + 6'b000101;
  assign Accum2_acc_1630_nl = nl_Accum2_acc_1630_nl[5:0];
  assign nl_Accum2_acc_1302_nl = conv_s2s_14_15(Product2_acc_792_cse_sva_1[15:2])
      + conv_s2s_13_15({Accum2_acc_1630_nl , (input_1_rsci_idat[58:52])}) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1);
  assign Accum2_acc_1302_nl = nl_Accum2_acc_1302_nl[14:0];
  assign nl_Accum2_acc_1304_nl = Product2_acc_1144_itm_16_1_1 + conv_s2s_15_16(Accum2_acc_1302_nl);
  assign Accum2_acc_1304_nl = nl_Accum2_acc_1304_nl[15:0];
  assign nl_Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1308_nl + Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_122_itm_17_2_1 + Accum2_acc_1305_nl + Accum2_acc_1304_nl + Product2_acc_367_itm_19_4_1
      + Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1 = (Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1631_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1[12:6])
      + 7'b0000001;
  assign Accum2_acc_1631_nl = nl_Accum2_acc_1631_nl[6:0];
  assign nl_Accum2_acc_1322_nl = conv_s2s_15_16(Product2_acc_609_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_1064_itm_16_1_1[15:1]) + conv_s2s_15_16(Product2_acc_33_itm_15_1_1)
      + conv_s2s_13_16({Accum2_acc_1631_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1[5:0])})
      + conv_s2s_13_16(input_1_rsci_idat[159:147]);
  assign Accum2_acc_1322_nl = nl_Accum2_acc_1322_nl[15:0];
  assign nl_Product2_acc_918_nl = conv_s2s_16_19(~ (input_1_rsci_idat[207:192]))
      + ({(input_1_rsci_idat[207:192]) , 3'b001});
  assign Product2_acc_918_nl = nl_Product2_acc_918_nl[18:0];
  assign nl_Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1322_nl + conv_s2s_14_16(Accum2_acc_1313_cse_1)
      + conv_s2s_14_16(input_1_rsci_idat[47:34]) + conv_s2s_15_16(readslicef_19_15_4(Product2_acc_918_nl))
      + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_934_itm_17_2_1[15:2]) + conv_s2s_14_16(Product2_acc_1334_itm_17_3_1[14:1]);
  assign Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1 = (Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product2_acc_1328_nl = conv_s2s_12_13(input_1_rsci_idat[159:148]) + 13'b0000000000001;
  assign Product2_acc_1328_nl = nl_Product2_acc_1328_nl[12:0];
  assign nl_Product2_acc_1280_nl = conv_s2s_16_17(input_1_rsci_idat[159:144]) + conv_s2s_15_17({Product2_acc_1328_nl
      , (input_1_rsci_idat[147:146])});
  assign Product2_acc_1280_nl = nl_Product2_acc_1280_nl[16:0];
  assign nl_Product2_acc_717_nl = conv_s2u_17_18(Product2_acc_1280_nl) + ({(~ (input_1_rsci_idat[159:144]))
      , 2'b00});
  assign Product2_acc_717_nl = nl_Product2_acc_717_nl[17:0];
  assign nl_Accum2_acc_1331_nl = Product2_acc_1084_itm_17_2_1 + (readslicef_18_16_2(Product2_acc_717_nl));
  assign Accum2_acc_1331_nl = nl_Accum2_acc_1331_nl[15:0];
  assign nl_Accum2_acc_1327_nl = conv_s2s_14_15(Product2_acc_943_cse_sva_1[15:2])
      + conv_s2s_13_15(input_1_rsci_idat[47:35]) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1);
  assign Accum2_acc_1327_nl = nl_Accum2_acc_1327_nl[14:0];
  assign nl_Accum2_acc_1330_nl = Product2_acc_1114_itm_17_2_1 + conv_s2s_15_16(Accum2_acc_1327_nl);
  assign Accum2_acc_1330_nl = nl_Accum2_acc_1330_nl[15:0];
  assign nl_Accum2_acc_1334_nl = Accum2_acc_1331_nl + Accum2_acc_1330_nl;
  assign Accum2_acc_1334_nl = nl_Accum2_acc_1334_nl[15:0];
  assign nl_Accum2_acc_1632_nl = conv_s2s_4_5(input_1_rsci_idat[143:140]) + 5'b00001;
  assign Accum2_acc_1632_nl = nl_Accum2_acc_1632_nl[4:0];
  assign nl_Accum2_acc_1333_nl = conv_s2s_15_16(Product2_acc_792_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_887_itm_15_1_1) + conv_s2s_15_16(Product2_acc_1332_itm_17_2_1[15:1])
      + conv_s2s_14_16(input_1_rsci_idat[15:2]) + conv_s2s_13_16({Accum2_acc_1632_nl
      , (input_1_rsci_idat[139:132])});
  assign Accum2_acc_1333_nl = nl_Accum2_acc_1333_nl[15:0];
  assign nl_Accum2_acc_1332_nl = Product2_acc_1053_itm_16_1_1 + Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1332_nl = nl_Accum2_acc_1332_nl[15:0];
  assign nl_Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1334_nl + Accum2_acc_1333_nl
      + Accum2_acc_1332_nl;
  assign Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1 = (Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1633_nl = conv_s2s_6_7(input_1_rsci_idat[207:202]) + 7'b1111001;
  assign Accum2_acc_1633_nl = nl_Accum2_acc_1633_nl[6:0];
  assign nl_Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_16(Product2_acc_478_itm_17_2_1[15:2]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(input_1_rsci_idat[47:33]) + conv_s2s_15_16(Product2_acc_1126_itm_16_1_1[15:1])
      + conv_s2s_13_16(Accum2_acc_1120_cse_1) + conv_s2s_13_16({Accum2_acc_1633_nl
      , (input_1_rsci_idat[201:196])}) + conv_s2s_13_16(input_1_rsci_idat[79:67])
      + conv_s2s_13_16(input_1_rsci_idat[127:115]);
  assign Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1 = (Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1354_nl = conv_s2s_15_16(Product2_acc_1126_itm_16_1_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_1334_itm_17_3_1) + conv_s2s_14_16(input_1_rsci_idat[79:66])
      + conv_s2s_14_16(Product2_acc_85_itm_15_1_1[14:1]);
  assign Accum2_acc_1354_nl = nl_Accum2_acc_1354_nl[15:0];
  assign nl_Accum2_acc_1353_nl = Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_216_itm_18_3_1[15:1]) + conv_s2s_15_16(Product2_acc_1042_itm_16_1_1[15:1]);
  assign Accum2_acc_1353_nl = nl_Accum2_acc_1353_nl[15:0];
  assign nl_Accum2_acc_1352_nl = Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_1118_itm_16_1_1;
  assign Accum2_acc_1352_nl = nl_Accum2_acc_1352_nl[15:0];
  assign nl_Accum2_acc_1351_nl = Product2_acc_954_itm_19_4_1 + conv_s2s_14_16(Product2_acc_867_cse_sva_1[15:2])
      + conv_s2s_14_16(Product2_acc_629_itm_17_3_1[14:1]);
  assign Accum2_acc_1351_nl = nl_Accum2_acc_1351_nl[15:0];
  assign nl_Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1354_nl + Accum2_acc_1353_nl
      + Accum2_acc_1352_nl + Accum2_acc_1351_nl;
  assign Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1 = (Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1366_nl = Accum2_acc_399_cse_1 + conv_s2s_15_16(input_1_rsci_idat[175:161])
      + conv_s2s_15_16(Product2_acc_1105_itm_16_1_1[15:1]);
  assign Accum2_acc_1366_nl = nl_Accum2_acc_1366_nl[15:0];
  assign nl_Accum2_acc_1365_nl = Product2_acc_152_itm_17_2_1 + Product2_acc_554_itm_19_4_1;
  assign Accum2_acc_1365_nl = nl_Accum2_acc_1365_nl[15:0];
  assign nl_Accum2_acc_1359_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(input_1_rsci_idat[79:67]);
  assign Accum2_acc_1359_nl = nl_Accum2_acc_1359_nl[13:0];
  assign nl_Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1366_nl + Accum2_acc_1365_nl
      + conv_s2s_14_16(Accum2_acc_1359_nl) + conv_s2s_14_16(input_1_rsci_idat[191:178])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[95:83]) + conv_s2s_13_16(input_1_rsci_idat[207:195]);
  assign Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1 = (Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1369_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[127:116]);
  assign Accum2_acc_1369_nl = nl_Accum2_acc_1369_nl[12:0];
  assign nl_Accum2_acc_1378_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_195_cse_sva_1[15:1]) + conv_s2s_15_16(Product2_acc_itm_18_3_1[15:1])
      + conv_s2s_14_16(Product2_acc_122_itm_17_2_1[15:2]) + conv_s2s_13_16(Accum2_acc_1369_nl);
  assign Accum2_acc_1378_nl = nl_Accum2_acc_1378_nl[15:0];
  assign nl_Accum2_acc_1634_nl = conv_s2s_4_5(input_1_rsci_idat[175:172]) + 5'b11111;
  assign Accum2_acc_1634_nl = nl_Accum2_acc_1634_nl[4:0];
  assign nl_Accum2_acc_1373_nl = (Product2_acc_1034_itm_16_1_1[15:1]) + conv_s2s_13_15({Accum2_acc_1634_nl
      , (input_1_rsci_idat[171:164])}) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1);
  assign Accum2_acc_1373_nl = nl_Accum2_acc_1373_nl[14:0];
  assign nl_Accum2_acc_1377_nl = conv_s2s_15_16(Accum2_acc_1373_nl) + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1377_nl = nl_Accum2_acc_1377_nl[15:0];
  assign nl_Accum2_acc_1376_nl = Product2_acc_367_itm_19_4_1 + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_447_itm_15_1_1[14:1]);
  assign Accum2_acc_1376_nl = nl_Accum2_acc_1376_nl[15:0];
  assign nl_Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1378_nl + Accum2_acc_1377_nl
      + Accum2_acc_1376_nl;
  assign Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1 = (Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1635_nl = conv_s2s_6_7(input_1_rsci_idat[95:90]) + 7'b0000101;
  assign Accum2_acc_1635_nl = nl_Accum2_acc_1635_nl[6:0];
  assign nl_Accum2_acc_1382_nl = conv_s2s_14_15(Product2_acc_730_cse_sva_1[15:2])
      + conv_s2s_13_15({Accum2_acc_1635_nl , (input_1_rsci_idat[89:84])}) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1);
  assign Accum2_acc_1382_nl = nl_Accum2_acc_1382_nl[14:0];
  assign nl_Accum2_acc_1385_nl = Product2_acc_943_cse_sva_1 + conv_s2s_15_16(Accum2_acc_1382_nl);
  assign Accum2_acc_1385_nl = nl_Accum2_acc_1385_nl[15:0];
  assign nl_Accum2_acc_1389_nl = Accum2_acc_1385_nl + conv_s2s_15_16(Product2_acc_667_cse_sva_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1389_nl = nl_Accum2_acc_1389_nl[15:0];
  assign Product2_acc_1329_nl =  -conv_s2s_14_15(input_1_rsci_idat[47:34]);
  assign nl_Product2_acc_182_nl = conv_s2s_17_19({Product2_acc_1329_nl , (~ (input_1_rsci_idat[33:32]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[47:32])) , 2'b01});
  assign Product2_acc_182_nl = nl_Product2_acc_182_nl[18:0];
  assign nl_Accum2_acc_1388_nl = (readslicef_19_16_3(Product2_acc_182_nl)) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_3_itm_15_1_1);
  assign Accum2_acc_1388_nl = nl_Accum2_acc_1388_nl[15:0];
  assign nl_Accum2_acc_1387_nl = Product2_acc_238_itm_17_2_1 + Product2_acc_455_itm_19_4_1;
  assign Accum2_acc_1387_nl = nl_Accum2_acc_1387_nl[15:0];
  assign nl_Product2_acc_1282_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[207:192]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[207:192]));
  assign Product2_acc_1282_nl = nl_Product2_acc_1282_nl[18:0];
  assign nl_Product2_acc_922_nl = conv_s2s_19_20(Product2_acc_1282_nl) + ({(input_1_rsci_idat[207:192])
      , 4'b0100});
  assign Product2_acc_922_nl = nl_Product2_acc_922_nl[19:0];
  assign nl_Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1389_nl + Accum2_acc_1388_nl
      + Accum2_acc_1387_nl + Product2_acc_834_itm_19_4_1 + (readslicef_20_16_4(Product2_acc_922_nl));
  assign Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1 = (Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1399_nl = Product2_acc_367_itm_19_4_1 + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_204_cse_sva_1[15:1]);
  assign Accum2_acc_1399_nl = nl_Accum2_acc_1399_nl[15:0];
  assign nl_Accum2_acc_1636_nl = conv_s2s_6_7(input_1_rsci_idat[79:74]) + 7'b0001101;
  assign Accum2_acc_1636_nl = nl_Accum2_acc_1636_nl[6:0];
  assign nl_Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1399_nl + Product2_acc_769_itm_19_4_1
      + Product2_acc_952_itm_19_4_1 + Product2_acc_458_itm_18_3_1 + Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_15_16(Product2_acc_887_itm_15_1_1) + conv_s2s_14_16(input_1_rsci_idat[47:34])
      + conv_s2s_13_16({Accum2_acc_1636_nl , (input_1_rsci_idat[73:68])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1 = (Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1412_nl = conv_s2s_15_16(Product2_acc_796_itm_18_4_1) + conv_s2s_15_16(Product2_acc_733_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_1147_itm_16_2_1) + conv_s2s_14_16(Product2_acc_308_cse_sva_1[15:2])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1);
  assign Accum2_acc_1412_nl = nl_Accum2_acc_1412_nl[15:0];
  assign nl_Accum2_acc_1404_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_129_12_8 , (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[7:0])});
  assign Accum2_acc_1404_nl = nl_Accum2_acc_1404_nl[13:0];
  assign nl_Accum2_acc_1411_nl = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(input_1_rsci_idat[15:1]) + conv_s2s_14_16(Accum2_acc_1404_nl);
  assign Accum2_acc_1411_nl = nl_Accum2_acc_1411_nl[15:0];
  assign nl_Accum2_acc_1410_nl = Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_1101_itm_16_1_1;
  assign Accum2_acc_1410_nl = nl_Accum2_acc_1410_nl[15:0];
  assign nl_Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1412_nl + Accum2_acc_1411_nl
      + Accum2_acc_1410_nl;
  assign Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1539_nl = conv_s2s_6_7(input_1_rsci_idat[143:138]) + 7'b0000001;
  assign Accum2_acc_1539_nl = nl_Accum2_acc_1539_nl[6:0];
  assign nl_Accum2_acc_nl = conv_s2s_15_16(Product2_acc_666_itm_18_3_1[15:1]) + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(Product2_acc_85_itm_15_1_1) + conv_s2s_13_16({Accum2_acc_1539_nl
      , (input_1_rsci_idat[137:132])}) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1);
  assign Accum2_acc_nl = nl_Accum2_acc_nl[15:0];
  assign nl_Accum2_acc_204_nl = conv_s2s_14_15(input_1_rsci_idat[207:194]) + conv_s2s_14_15(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_204_nl = nl_Accum2_acc_204_nl[14:0];
  assign nl_Accum2_acc_208_nl = Product2_acc_492_itm_17_2_1 + conv_s2s_15_16(Accum2_acc_204_nl);
  assign Accum2_acc_208_nl = nl_Accum2_acc_208_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1 = Accum2_acc_nl
      + Accum2_acc_208_nl + conv_s2s_15_16(input_1_rsci_idat[63:49]) + conv_s2s_14_16(Product2_acc_370_cse_sva_1[15:2])
      + conv_s2s_14_16(Product2_acc_1338_itm_17_3_1[14:1]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1 = (Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1424_nl = Accum2_acc_1066_cse_1 + conv_s2s_15_16(input_1_rsci_idat[127:113])
      + conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1]);
  assign Accum2_acc_1424_nl = nl_Accum2_acc_1424_nl[15:0];
  assign nl_Accum2_acc_1638_nl = conv_s2s_6_7(input_1_rsci_idat[143:138]) + 7'b0000011;
  assign Accum2_acc_1638_nl = nl_Accum2_acc_1638_nl[6:0];
  assign nl_Accum2_acc_1415_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1638_nl , (input_1_rsci_idat[137:132])});
  assign Accum2_acc_1415_nl = nl_Accum2_acc_1415_nl[13:0];
  assign nl_Accum2_acc_1423_nl = conv_s2s_15_16(Product2_acc_728_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_797_cse_sva_1[15:1]) + conv_s2s_15_16(Product2_acc_3_itm_15_1_1)
      + conv_s2s_14_16(Accum2_acc_1415_nl);
  assign Accum2_acc_1423_nl = nl_Accum2_acc_1423_nl[15:0];
  assign nl_Accum2_acc_1416_nl = conv_s2s_14_15(input_1_rsci_idat[47:34]) + conv_s2s_14_15(Product2_acc_1330_itm_17_3_1[14:1]);
  assign Accum2_acc_1416_nl = nl_Accum2_acc_1416_nl[14:0];
  assign nl_Accum2_acc_1421_nl = Product2_acc_1144_itm_16_1_1 + conv_s2s_15_16(Accum2_acc_1416_nl);
  assign Accum2_acc_1421_nl = nl_Accum2_acc_1421_nl[15:0];
  assign nl_Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1424_nl + Accum2_acc_1423_nl
      + Accum2_acc_1421_nl + Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_283_itm_18_3_1;
  assign Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1 = (Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1433_nl = Product2_acc_1117_itm_16_1_1 + Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1433_nl = nl_Accum2_acc_1433_nl[15:0];
  assign nl_Accum2_acc_1437_nl = Accum2_acc_1433_nl + conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1])
      + conv_s2s_14_16(input_1_rsci_idat[143:130]) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1437_nl = nl_Accum2_acc_1437_nl[15:0];
  assign nl_Accum2_acc_1639_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1[12:7])
      + 6'b000001;
  assign Accum2_acc_1639_nl = nl_Accum2_acc_1639_nl[5:0];
  assign nl_Accum2_acc_1436_nl = conv_s2s_15_16(Product2_acc_796_itm_18_4_1) + conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_195_cse_sva_1[15:1]) + conv_s2s_13_16({Accum2_acc_1639_nl
      , (nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1[6:0])})
      + conv_s2s_13_16(input_1_rsci_idat[15:3]);
  assign Accum2_acc_1436_nl = nl_Accum2_acc_1436_nl[15:0];
  assign nl_Accum2_acc_1434_nl = Product2_acc_532_cse_sva_1 + Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1434_nl = nl_Accum2_acc_1434_nl[15:0];
  assign nl_Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1437_nl + Accum2_acc_1436_nl
      + Accum2_acc_1434_nl + Product2_acc_297_itm_17_2_1 + Product2_acc_476_itm_19_4_1;
  assign Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1 = (Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1446_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_14_15(Accum2_acc_1028_cse_1);
  assign Accum2_acc_1446_nl = nl_Accum2_acc_1446_nl[14:0];
  assign nl_Accum2_acc_1448_nl = Product2_acc_531_itm_19_4_1 + conv_s2s_15_16(Accum2_acc_1446_nl);
  assign Accum2_acc_1448_nl = nl_Accum2_acc_1448_nl[15:0];
  assign nl_Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1448_nl + Product2_acc_299_itm_19_4_1
      + Product2_acc_450_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_476_cse_1) + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1)
      + conv_s2s_13_16(input_1_rsci_idat[175:163]);
  assign Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1 = (Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1460_nl = conv_s2s_15_16(input_1_rsci_idat[159:145]) + conv_s2s_15_16(Product2_acc_216_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_1027_itm_16_2_1) + conv_s2s_14_16(Product2_acc_733_itm_17_2_1[15:2])
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1460_nl = nl_Accum2_acc_1460_nl[15:0];
  assign nl_Accum2_acc_1459_nl = Product2_acc_1034_itm_16_1_1 + Product2_acc_285_itm_19_4_1;
  assign Accum2_acc_1459_nl = nl_Accum2_acc_1459_nl[15:0];
  assign nl_Accum2_acc_1458_nl = Product2_acc_368_cse_sva_1 + Product2_acc_478_itm_17_2_1;
  assign Accum2_acc_1458_nl = nl_Accum2_acc_1458_nl[15:0];
  assign nl_Accum2_acc_1457_nl = Product2_acc_946_itm_18_3_1 + conv_s2s_14_16(input_1_rsci_idat[127:114])
      + conv_s2s_13_16({Accum2_Accum2_conc_111_12_7 , (input_1_rsci_idat[186:180])})
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1);
  assign Accum2_acc_1457_nl = nl_Accum2_acc_1457_nl[15:0];
  assign nl_Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1460_nl + Accum2_acc_1459_nl
      + Accum2_acc_1458_nl + Accum2_acc_1457_nl;
  assign Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1 = (Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1471_nl = Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_532_cse_sva_1;
  assign Accum2_acc_1471_nl = nl_Accum2_acc_1471_nl[15:0];
  assign nl_Accum2_acc_1470_nl = Product2_acc_792_cse_sva_1 + Product2_acc_1144_itm_16_1_1;
  assign Accum2_acc_1470_nl = nl_Accum2_acc_1470_nl[15:0];
  assign nl_Accum2_acc_1474_nl = Accum2_acc_1471_nl + Accum2_acc_1470_nl;
  assign Accum2_acc_1474_nl = nl_Accum2_acc_1474_nl[15:0];
  assign nl_Accum2_acc_1642_nl = conv_s2s_4_5(input_1_rsci_idat[31:28]) + 5'b00001;
  assign Accum2_acc_1642_nl = nl_Accum2_acc_1642_nl[4:0];
  assign nl_Accum2_acc_1473_nl = conv_s2s_15_16(input_1_rsci_idat[15:1]) + conv_s2s_15_16(input_1_rsci_idat[95:81])
      + conv_s2s_14_16(input_1_rsci_idat[143:130]) + conv_s2s_14_16(Product2_acc_871_itm_17_2_1[15:2])
      + conv_s2s_14_16(Product2_acc_122_itm_17_2_1[15:2]) + conv_s2s_13_16({Accum2_acc_1642_nl
      , (input_1_rsci_idat[27:20])});
  assign Accum2_acc_1473_nl = nl_Accum2_acc_1473_nl[15:0];
  assign nl_Accum2_acc_1467_nl = conv_s2s_15_16(Product2_acc_1064_itm_16_1_1[15:1])
      + conv_s2s_13_16(input_1_rsci_idat[175:163]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1);
  assign Accum2_acc_1467_nl = nl_Accum2_acc_1467_nl[15:0];
  assign nl_Accum2_acc_1472_nl = Accum2_acc_1467_nl + Product2_acc_1056_itm_16_1_1;
  assign Accum2_acc_1472_nl = nl_Accum2_acc_1472_nl[15:0];
  assign nl_Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1474_nl + Accum2_acc_1473_nl
      + Accum2_acc_1472_nl;
  assign Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1 = (Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_249_nl = conv_s2s_12_13(input_1_rsci_idat[143:132])
      + 13'b0000110000001;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_249_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_249_nl[12:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_257_nl = Product2_acc_952_itm_19_4_1
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_249_nl)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_257_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_257_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_260_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_257_nl
      + conv_s2s_15_16(Product2_acc_802_itm_17_2_1[15:1]) + conv_s2s_15_16(Product2_acc_290_itm_15_1_1);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_260_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_260_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_251_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[15:4]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_251_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_251_nl[12:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_255_nl = conv_s2s_15_16(Product2_acc_217_itm_17_2_1[15:1])
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_251_nl)
      + conv_s2s_12_16(input_1_rsci_idat[47:36]) + conv_s2s_12_16(input_1_rsci_idat[127:116]);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_255_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_255_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_259_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_255_nl
      + (~ (input_1_rsci_idat[175:160]));
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_259_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_259_nl[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_258_nl = Product2_acc_1080_itm_16_1_1
      + Product2_acc_691_itm_19_4_1;
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_258_nl = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_258_nl[15:0];
  assign nl_Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_260_nl
      + nnet_product_mult_input_t_config2_weight_t_product_acc_259_nl + nnet_product_mult_input_t_config2_weight_t_product_acc_258_nl;
  assign Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1 = (Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1643_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[12:7])
      + 6'b111001;
  assign Accum2_acc_1643_nl = nl_Accum2_acc_1643_nl[5:0];
  assign nl_Accum1_2_Accum2_123_Accum2_acc_1_nl = conv_s2s_13_15({Accum2_acc_1643_nl
      , (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[6:0])})
      + Product2_acc_1027_itm_16_2_1;
  assign Accum1_2_Accum2_123_Accum2_acc_1_nl = nl_Accum1_2_Accum2_123_Accum2_acc_1_nl[14:0];
  assign nl_Accum2_acc_1481_nl = conv_s2s_15_16(Product2_acc_124_cse_sva_1[15:1])
      + conv_s2s_15_16(Accum1_2_Accum2_123_Accum2_acc_1_nl);
  assign Accum2_acc_1481_nl = nl_Accum2_acc_1481_nl[15:0];
  assign nl_Accum2_acc_1483_nl = Accum2_acc_1481_nl + Product2_acc_195_cse_sva_1;
  assign Accum2_acc_1483_nl = nl_Accum2_acc_1483_nl[15:0];
  assign nl_Accum2_acc_1477_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[95:84]);
  assign Accum2_acc_1477_nl = nl_Accum2_acc_1477_nl[12:0];
  assign nl_Accum2_acc_1479_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14(Accum2_acc_1477_nl);
  assign Accum2_acc_1479_nl = nl_Accum2_acc_1479_nl[13:0];
  assign nl_Accum2_acc_1480_nl = conv_s2s_14_15(Accum2_acc_1479_nl) + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1)
      + conv_s2s_13_15(nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1);
  assign Accum2_acc_1480_nl = nl_Accum2_acc_1480_nl[14:0];
  assign nl_Accum2_acc_1482_nl = Product2_acc_308_cse_sva_1 + conv_s2s_15_16(Accum2_acc_1480_nl);
  assign Accum2_acc_1482_nl = nl_Accum2_acc_1482_nl[15:0];
  assign nl_Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1483_nl + Accum2_acc_1482_nl;
  assign Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1 = (Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1644_nl = (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[12:6])
      + 7'b0000101;
  assign Accum2_acc_1644_nl = nl_Accum2_acc_1644_nl[6:0];
  assign nl_Accum2_acc_1492_nl = conv_s2s_15_16(Product2_acc_1086_itm_16_1_1[15:1])
      + conv_s2s_15_16(Product2_acc_1042_itm_16_1_1[15:1]) + conv_s2s_14_16(input_1_rsci_idat[207:194])
      + conv_s2s_13_16({Accum2_acc_1644_nl , (nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[5:0])})
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1)
      + conv_s2s_14_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_377_itm_17_2_1[15:2]);
  assign Accum2_acc_1492_nl = nl_Accum2_acc_1492_nl[15:0];
  assign nl_Accum2_acc_1491_nl = Product2_acc_75_itm_19_4_1 + Product2_acc_1056_itm_16_1_1;
  assign Accum2_acc_1491_nl = nl_Accum2_acc_1491_nl[15:0];
  assign nl_Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1492_nl + Accum2_acc_1491_nl
      + Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_946_itm_18_3_1;
  assign Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1 = (Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1645_nl = conv_s2s_6_7(input_1_rsci_idat[207:202]) + 7'b1111011;
  assign Accum2_acc_1645_nl = nl_Accum2_acc_1645_nl[6:0];
  assign nl_Accum2_acc_1496_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_acc_1645_nl , (input_1_rsci_idat[201:196])});
  assign Accum2_acc_1496_nl = nl_Accum2_acc_1496_nl[13:0];
  assign nl_Accum2_acc_1501_nl = Product2_acc_834_itm_19_4_1 + conv_s2s_14_16(Accum2_acc_1496_nl)
      + conv_s2s_13_16(input_1_rsci_idat[127:115]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1);
  assign Accum2_acc_1501_nl = nl_Accum2_acc_1501_nl[15:0];
  assign nl_Accum2_acc_1504_nl = Accum2_acc_1501_nl + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(input_1_rsci_idat[63:50]) + conv_s2s_14_16(Product2_acc_934_itm_17_2_1[15:2]);
  assign Accum2_acc_1504_nl = nl_Accum2_acc_1504_nl[15:0];
  assign nl_Accum2_acc_1503_nl = Product2_acc_75_itm_19_4_1 + conv_s2s_15_16(Product2_acc_297_itm_17_2_1[15:1])
      + conv_s2s_15_16(Product2_acc_33_itm_15_1_1);
  assign Accum2_acc_1503_nl = nl_Accum2_acc_1503_nl[15:0];
  assign nl_Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1504_nl + Accum2_acc_1503_nl
      + Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_728_itm_18_3_1;
  assign Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1 = (Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1514_nl = Product2_acc_1034_itm_16_1_1 + Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1;
  assign Accum2_acc_1514_nl = nl_Accum2_acc_1514_nl[15:0];
  assign nl_Accum2_acc_1507_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[47:36]);
  assign Accum2_acc_1507_nl = nl_Accum2_acc_1507_nl[12:0];
  assign nl_Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1514_nl + conv_s2s_15_16(Product2_acc_478_itm_17_2_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_14_16(Product2_acc_195_cse_sva_1[15:2]) + conv_s2s_13_16(Accum2_acc_1507_nl)
      + conv_s2s_13_16({Accum2_Accum2_conc_125_12_6 , (input_1_rsci_idat[217:212])})
      + conv_s2s_13_16(input_1_rsci_idat[127:115]) + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1)
      + conv_s2s_13_16(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1);
  assign Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1 = (Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1517_nl = nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[47:36]);
  assign Accum2_acc_1517_nl = nl_Accum2_acc_1517_nl[12:0];
  assign nl_Accum2_acc_1525_nl = Accum2_acc_411_cse_1 + conv_s2s_15_16(Product2_acc_308_cse_sva_1[15:1])
      + conv_s2s_13_16(Accum2_acc_1517_nl) + conv_s2s_13_16({Accum2_Accum2_conc_125_12_6
      , (input_1_rsci_idat[217:212])});
  assign Accum2_acc_1525_nl = nl_Accum2_acc_1525_nl[15:0];
  assign nl_Accum2_acc_1524_nl = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + Product2_acc_532_cse_sva_1;
  assign Accum2_acc_1524_nl = nl_Accum2_acc_1524_nl[15:0];
  assign nl_Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1525_nl + Accum2_acc_1524_nl
      + conv_s2s_15_16(Product2_acc_1134_itm_16_1_1[15:1]) + conv_s2s_14_16(Accum2_acc_1313_cse_1)
      + conv_s2s_14_16(Product2_acc_478_itm_17_2_1[15:2]);
  assign Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 = (Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Accum2_acc_1537_nl = conv_s2s_15_16(Product2_acc_1110_itm_16_2_1) + conv_s2s_15_16(Product2_acc_1064_itm_16_1_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_1537_nl = nl_Accum2_acc_1537_nl[15:0];
  assign nl_Accum1_2_Accum2_128_Accum2_acc_1_nl = conv_s2s_14_15({Accum2_acc_1558_cse_1
      , (input_1_rsci_idat[25:19])}) + Product2_acc_1027_itm_16_2_1;
  assign Accum1_2_Accum2_128_Accum2_acc_1_nl = nl_Accum1_2_Accum2_128_Accum2_acc_1_nl[14:0];
  assign nl_Accum2_acc_1536_nl = conv_s2s_15_16(Accum1_2_Accum2_128_Accum2_acc_1_nl)
      + conv_s2s_14_16(input_1_rsci_idat[175:162]) + conv_s2s_14_16(Product2_acc_792_cse_sva_1[15:2])
      + conv_s2s_13_16(input_1_rsci_idat[207:195]) + conv_s2s_12_16(input_1_rsci_idat[127:116])
      + conv_s2s_12_16(input_1_rsci_idat[143:132]);
  assign Accum2_acc_1536_nl = nl_Accum2_acc_1536_nl[15:0];
  assign nl_Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1537_nl + Accum2_acc_1536_nl
      + conv_s2s_15_16(Product2_acc_946_itm_18_3_1[15:1]) + conv_s2s_14_16(Product2_acc_478_itm_17_2_1[15:2])
      + conv_s2s_14_16(Product2_acc_377_itm_17_2_1[15:2]);
  assign Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_415_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_415_nl = nl_Product2_1_acc_415_nl[13:0];
  assign Product2_1_acc_415_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_415_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_418_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_418_nl = nl_Product2_1_acc_418_nl[12:0];
  assign Product2_1_acc_418_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_418_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_722_cse_1 = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_722_cse_1 = nl_Product2_1_acc_722_cse_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_423_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_423_nl = nl_Product2_1_acc_423_nl[12:0];
  assign Product2_1_acc_423_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_423_nl);
  assign nl_Product2_1_acc_424_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_424_nl = nl_Product2_1_acc_424_nl[13:0];
  assign Product2_1_acc_424_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_424_nl);
  assign nl_Product2_1_acc_425_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_425_nl = nl_Product2_1_acc_425_nl[13:0];
  assign Product2_1_acc_425_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_425_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_428_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_428_nl = nl_Product2_1_acc_428_nl[12:0];
  assign Product2_1_acc_428_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_428_nl);
  assign nl_Product2_1_acc_429_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_429_nl = nl_Product2_1_acc_429_nl[12:0];
  assign Product2_1_acc_429_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_429_nl);
  assign nl_Product2_1_acc_430_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_430_nl = nl_Product2_1_acc_430_nl[13:0];
  assign Product2_1_acc_430_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_430_nl);
  assign nl_Product2_1_acc_431_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_431_nl = nl_Product2_1_acc_431_nl[12:0];
  assign Product2_1_acc_431_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_431_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_67_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_67_nl = nl_Product2_1_acc_67_nl[11:0];
  assign Product2_1_acc_67_itm_11_4_1 = readslicef_12_8_4(Product2_1_acc_67_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_384_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_384_nl = nl_Product2_1_acc_384_nl[10:0];
  assign Product2_1_acc_384_itm_10_1_1 = readslicef_11_10_1(Product2_1_acc_384_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_396_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_396_nl = nl_Product2_1_acc_396_nl[12:0];
  assign Product2_1_acc_396_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_396_nl);
  assign nl_Product2_1_acc_76_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_76_nl = nl_Product2_1_acc_76_nl[11:0];
  assign Product2_1_acc_76_itm_11_4_1 = readslicef_12_8_4(Product2_1_acc_76_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_391_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_391_nl = nl_Product2_1_acc_391_nl[12:0];
  assign Product2_1_acc_391_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_391_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_393_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_393_nl = nl_Product2_1_acc_393_nl[12:0];
  assign Product2_1_acc_393_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_393_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_399_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_399_nl = nl_Product2_1_acc_399_nl[12:0];
  assign Product2_1_acc_399_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_399_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_478_nl = conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_478_nl = nl_Product2_1_acc_478_nl[10:0];
  assign Product2_1_acc_478_itm_10_2_1 = readslicef_11_9_2(Product2_1_acc_478_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_72_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_72_nl = nl_Product2_1_acc_72_nl[11:0];
  assign Product2_1_acc_72_itm_11_3_1 = readslicef_12_9_3(Product2_1_acc_72_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_241_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_241_nl = nl_Product2_1_acc_241_nl[11:0];
  assign Product2_1_acc_241_itm_11_4_1 = readslicef_12_8_4(Product2_1_acc_241_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1);
  assign layer4_out_0_9_1_lpi_1_dfm_1 = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_0_0_lpi_1_dfm_1 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_469_nl = conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_469_nl = nl_Product2_1_acc_469_nl[10:0];
  assign Product2_1_acc_469_itm_10_1_1 = readslicef_11_10_1(Product2_1_acc_469_nl);
  assign nl_Product2_1_acc_8_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_8_nl = nl_Product2_1_acc_8_nl[11:0];
  assign Product2_1_acc_8_itm_11_2_1 = readslicef_12_10_2(Product2_1_acc_8_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      = (Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1
      = MUX_v_9_2_2(9'b000000000, ({nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_nl
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl}),
      nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_410_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_410_nl = nl_Product2_1_acc_410_nl[13:0];
  assign Product2_1_acc_410_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_410_nl);
  assign nl_Product2_1_acc_411_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_411_nl = nl_Product2_1_acc_411_nl[13:0];
  assign Product2_1_acc_411_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_411_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_414_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_414_nl = nl_Product2_1_acc_414_nl[12:0];
  assign Product2_1_acc_414_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_414_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_9
      = ((Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_0
      = ((Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_644_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_949 , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_949});
  assign Product2_1_acc_644_nl = nl_Product2_1_acc_644_nl[13:0];
  assign Product2_1_acc_644_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_644_nl);
  assign nl_Product2_1_acc_645_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_943 , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_943});
  assign Product2_1_acc_645_nl = nl_Product2_1_acc_645_nl[12:0];
  assign Product2_1_acc_645_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_645_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_633_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_633_nl = nl_Product2_1_acc_633_nl[12:0];
  assign Product2_1_acc_633_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_633_nl);
  assign nl_Product2_1_acc_634_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_634_nl = nl_Product2_1_acc_634_nl[12:0];
  assign Product2_1_acc_634_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_634_nl);
  assign nl_Product2_1_acc_636_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_636_nl = nl_Product2_1_acc_636_nl[12:0];
  assign Product2_1_acc_636_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_636_nl);
  assign nl_Product2_1_acc_638_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_638_nl = nl_Product2_1_acc_638_nl[12:0];
  assign Product2_1_acc_638_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_638_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_641_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_941 , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_941});
  assign Product2_1_acc_641_nl = nl_Product2_1_acc_641_nl[12:0];
  assign Product2_1_acc_641_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_641_nl);
  assign nl_Product2_1_acc_642_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_642_nl = nl_Product2_1_acc_642_nl[12:0];
  assign Product2_1_acc_642_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_642_nl);
  assign nl_Product2_1_acc_79_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_79_nl = nl_Product2_1_acc_79_nl[11:0];
  assign Product2_1_acc_79_itm_11_4_1 = readslicef_12_8_4(Product2_1_acc_79_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_41_nl = ~((((Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1)
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1
      = ({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2s_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_41_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1[7:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_25_nl = ~((((nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1)
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1
      = ({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2s_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_25_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_643_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_643_nl = nl_Product2_1_acc_643_nl[13:0];
  assign Product2_1_acc_643_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_643_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_476_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_476_nl = nl_Product2_1_acc_476_nl[13:0];
  assign Product2_1_acc_476_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_476_nl);
  assign nl_Product2_1_acc_477_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_963 , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_963});
  assign Product2_1_acc_477_nl = nl_Product2_1_acc_477_nl[13:0];
  assign Product2_1_acc_477_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_477_nl);
  assign nl_Product2_1_acc_480_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_480_nl = nl_Product2_1_acc_480_nl[13:0];
  assign Product2_1_acc_480_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_480_nl);
  assign nl_Product2_1_acc_483_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_483_nl = nl_Product2_1_acc_483_nl[13:0];
  assign Product2_1_acc_483_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_483_nl);
  assign nl_Product2_1_acc_484_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_484_nl = nl_Product2_1_acc_484_nl[12:0];
  assign Product2_1_acc_484_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_484_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_450_nl = conv_u2u_12_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_not_279
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_not_279
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_450_nl = nl_Product2_1_acc_450_nl[12:0];
  assign Product2_1_acc_450_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_450_nl);
  assign nl_Product2_1_acc_462_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_462_nl = nl_Product2_1_acc_462_nl[12:0];
  assign Product2_1_acc_462_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_462_nl);
  assign nl_Product2_1_acc_464_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_464_nl = nl_Product2_1_acc_464_nl[12:0];
  assign Product2_1_acc_464_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_464_nl);
  assign nl_Product2_1_acc_454_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_454_nl = nl_Product2_1_acc_454_nl[12:0];
  assign Product2_1_acc_454_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_454_nl);
  assign nl_Product2_1_acc_455_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_911 , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_911});
  assign Product2_1_acc_455_nl = nl_Product2_1_acc_455_nl[12:0];
  assign Product2_1_acc_455_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_455_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nl_Product2_1_acc_466_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_466_nl = nl_Product2_1_acc_466_nl[13:0];
  assign Product2_1_acc_466_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_466_nl);
  assign nl_Product2_1_acc_467_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_467_nl = nl_Product2_1_acc_467_nl[12:0];
  assign Product2_1_acc_467_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_467_nl);
  assign nl_Product2_1_acc_468_nl = conv_u2u_13_14({(~ layer4_out_0_9_1_lpi_1_dfm_1)
      , (~ layer4_out_0_0_lpi_1_dfm_1) , 3'b001}) + conv_u2u_10_14({(~ layer4_out_0_9_1_lpi_1_dfm_1)
      , (~ layer4_out_0_0_lpi_1_dfm_1)});
  assign Product2_1_acc_468_nl = nl_Product2_1_acc_468_nl[13:0];
  assign Product2_1_acc_468_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_468_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nl_Product2_1_acc_473_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_473_nl = nl_Product2_1_acc_473_nl[13:0];
  assign Product2_1_acc_473_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_473_nl);
  assign nl_Product2_1_acc_474_nl = conv_u2u_13_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 3'b001}) + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_474_nl = nl_Product2_1_acc_474_nl[13:0];
  assign Product2_1_acc_474_itm_13_3_1 = readslicef_14_11_3(Product2_1_acc_474_nl);
  assign nl_Product2_1_acc_475_nl = conv_u2u_12_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b01}) + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_475_nl = nl_Product2_1_acc_475_nl[12:0];
  assign Product2_1_acc_475_itm_12_2_1 = readslicef_13_11_2(Product2_1_acc_475_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_9_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_8_1_lpi_1_dfm_1
      = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_1_pmx_0_lpi_1_dfm_1
      = ((nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_115_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nl_Accum2_acc_1558_cse_1 = conv_s2u_6_7(input_1_rsci_idat[31:26]) + 7'b1111011;
  assign Accum2_acc_1558_cse_1 = nl_Accum2_acc_1558_cse_1[6:0];
  assign nl_Product2_acc_1027_nl = conv_s2u_14_17(input_1_rsci_idat[15:2]) + conv_s2u_16_17(input_1_rsci_idat[15:0]);
  assign Product2_acc_1027_nl = nl_Product2_acc_1027_nl[16:0];
  assign Product2_acc_1027_itm_16_2_1 = readslicef_17_15_2(Product2_acc_1027_nl);
  assign nl_Product2_acc_792_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[191:178])
      - (input_1_rsci_idat[191:176]);
  assign Product2_acc_792_cse_sva_1 = nl_Product2_acc_792_cse_sva_1[15:0];
  assign nl_Product2_acc_478_nl = conv_s2s_16_18(~ (input_1_rsci_idat[111:96])) +
      ({(input_1_rsci_idat[111:96]) , 2'b01});
  assign Product2_acc_478_nl = nl_Product2_acc_478_nl[17:0];
  assign Product2_acc_478_itm_17_2_1 = readslicef_18_16_2(Product2_acc_478_nl);
  assign nl_Product2_acc_377_nl = conv_s2s_16_18(~ (input_1_rsci_idat[95:80])) +
      ({(input_1_rsci_idat[95:80]) , 2'b01});
  assign Product2_acc_377_nl = nl_Product2_acc_377_nl[17:0];
  assign Product2_acc_377_itm_17_2_1 = readslicef_18_16_2(Product2_acc_377_nl);
  assign nl_Product2_acc_946_nl = conv_s2s_16_19(~ (input_1_rsci_idat[223:208]))
      + ({(input_1_rsci_idat[223:208]) , 3'b001});
  assign Product2_acc_946_nl = nl_Product2_acc_946_nl[18:0];
  assign Product2_acc_946_itm_18_3_1 = readslicef_19_16_3(Product2_acc_946_nl);
  assign nl_Product2_acc_1064_nl = conv_s2u_14_17(input_1_rsci_idat[79:66]) + conv_s2u_16_17(input_1_rsci_idat[79:64]);
  assign Product2_acc_1064_nl = nl_Product2_acc_1064_nl[16:0];
  assign Product2_acc_1064_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1064_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_208_nl = ~((input_1_rsci_idat[33:32]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[47:34])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_208_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_219_nl = ~((input_1_rsci_idat[49:48]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[63:50])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_219_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[95:81])) + conv_u2s_1_16(~ (input_1_rsci_idat[80]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Product2_acc_532_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[127:114])
      - (input_1_rsci_idat[127:112]);
  assign Product2_acc_532_cse_sva_1 = nl_Product2_acc_532_cse_sva_1[15:0];
  assign nl_Accum2_acc_1313_cse_1 = conv_s2s_13_14(input_1_rsci_idat[191:179]) +
      conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1);
  assign Accum2_acc_1313_cse_1 = nl_Accum2_acc_1313_cse_1[13:0];
  assign nl_Product2_acc_1134_nl = conv_s2u_14_17(input_1_rsci_idat[207:194]) + conv_s2u_16_17(input_1_rsci_idat[207:192]);
  assign Product2_acc_1134_nl = nl_Product2_acc_1134_nl[16:0];
  assign Product2_acc_1134_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1134_nl);
  assign nl_Accum2_acc_411_cse_1 = conv_s2s_15_16(Product2_acc_604_itm_18_3_1[15:1])
      + conv_s2s_15_16(Product2_acc_72_itm_18_3_1[15:1]);
  assign Accum2_acc_411_cse_1 = nl_Accum2_acc_411_cse_1[15:0];
  assign nl_Product2_acc_308_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[79:66])
      - (input_1_rsci_idat[79:64]);
  assign Product2_acc_308_cse_sva_1 = nl_Product2_acc_308_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_53_nl = ~((input_1_rsci_idat[51:48]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[63:52])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_53_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_52_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_85_nl = ~((input_1_rsci_idat[131:128]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[143:132])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_85_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_84_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_99_nl = ~((input_1_rsci_idat[147:144]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[159:148])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_99_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1[12:0];
  assign nl_Product2_acc_195_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[63:50])
      - (input_1_rsci_idat[63:48]);
  assign Product2_acc_195_cse_sva_1 = nl_Product2_acc_195_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_60_nl = ~((input_1_rsci_idat[83:80]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[95:84])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_60_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_59_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_167_nl = ~((input_1_rsci_idat[1:0]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[15:2])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_167_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_1034_nl = conv_s2u_14_17(input_1_rsci_idat[31:18]) + conv_s2u_16_17(input_1_rsci_idat[31:16]);
  assign Product2_acc_1034_nl = nl_Product2_acc_1034_nl[16:0];
  assign Product2_acc_1034_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1034_nl);
  assign nl_Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[79:64]);
  assign Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Product2_acc_297_nl = conv_s2s_16_18(~ (input_1_rsci_idat[79:64])) +
      ({(input_1_rsci_idat[79:64]) , 2'b01});
  assign Product2_acc_297_nl = nl_Product2_acc_297_nl[17:0];
  assign Product2_acc_297_itm_17_2_1 = readslicef_18_16_2(Product2_acc_297_nl);
  assign nl_Product2_acc_75_nl = conv_s2s_16_20(~ (input_1_rsci_idat[31:16])) + ({(input_1_rsci_idat[31:16])
      , 4'b0001});
  assign Product2_acc_75_nl = nl_Product2_acc_75_nl[19:0];
  assign Product2_acc_75_itm_19_4_1 = readslicef_20_16_4(Product2_acc_75_nl);
  assign nl_Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[95:80]);
  assign Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign Product2_acc_1307_nl =  -conv_s2s_14_15(input_1_rsci_idat[175:162]);
  assign nl_Product2_acc_728_nl = conv_s2s_17_19({Product2_acc_1307_nl , (~ (input_1_rsci_idat[161:160]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[175:160])) , 2'b01});
  assign Product2_acc_728_nl = nl_Product2_acc_728_nl[18:0];
  assign Product2_acc_728_itm_18_3_1 = readslicef_19_16_3(Product2_acc_728_nl);
  assign nl_Product2_acc_834_nl = conv_s2s_16_20(~ (input_1_rsci_idat[191:176]))
      + ({(input_1_rsci_idat[191:176]) , 4'b0001});
  assign Product2_acc_834_nl = nl_Product2_acc_834_nl[19:0];
  assign Product2_acc_834_itm_19_4_1 = readslicef_20_16_4(Product2_acc_834_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_274_nl = ~((input_1_rsci_idat[130:128]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[143:131])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_274_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_66_nl = ~((input_1_rsci_idat[99:96]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[111:100])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_66_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_65_cse_sva_1[12:0];
  assign nl_Product2_acc_934_nl = conv_s2s_16_18(~ (input_1_rsci_idat[223:208]))
      + ({(input_1_rsci_idat[223:208]) , 2'b01});
  assign Product2_acc_934_nl = nl_Product2_acc_934_nl[17:0];
  assign Product2_acc_934_itm_17_2_1 = readslicef_18_16_2(Product2_acc_934_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_287_nl = ~((input_1_rsci_idat[145:144]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[159:146])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_287_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_1056_nl = conv_s2u_13_17(input_1_rsci_idat[63:51]) + conv_s2u_16_17(input_1_rsci_idat[63:48]);
  assign Product2_acc_1056_nl = nl_Product2_acc_1056_nl[16:0];
  assign Product2_acc_1056_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1056_nl);
  assign nl_Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[143:128]);
  assign Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_1_nl = ~((input_1_rsci_idat[3:0]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1 = conv_s2s_12_13(~
      (input_1_rsci_idat[15:4])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_1_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_132_nl = ~((input_1_rsci_idat[179:176]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1
      = conv_s2s_12_13(~ (input_1_rsci_idat[191:180])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_132_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_301_nl = ~((input_1_rsci_idat[162:160]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[175:163])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_301_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Product2_acc_1086_nl = conv_s2u_14_17(input_1_rsci_idat[111:98]) + conv_s2u_16_17(input_1_rsci_idat[111:96]);
  assign Product2_acc_1086_nl = nl_Product2_acc_1086_nl[16:0];
  assign Product2_acc_1086_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1086_nl);
  assign nl_Product2_acc_1042_nl = conv_s2u_14_17(input_1_rsci_idat[47:34]) + conv_s2u_16_17(input_1_rsci_idat[47:32]);
  assign Product2_acc_1042_nl = nl_Product2_acc_1042_nl[16:0];
  assign Product2_acc_1042_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1042_nl);
  assign nl_Product2_acc_124_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[47:34])
      - (input_1_rsci_idat[47:32]);
  assign Product2_acc_124_cse_sva_1 = nl_Product2_acc_124_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_15_nl = ~((input_1_rsci_idat[19:16]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[31:20])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_15_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_336_nl = ~((input_1_rsci_idat[210:208]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[223:211])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_336_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_74_nl = ~((input_1_rsci_idat[115:112]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[127:116])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_74_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_121_nl = ~((input_1_rsci_idat[163:160]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1
      = conv_s2s_12_13(~ (input_1_rsci_idat[175:164])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_121_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1[12:0];
  assign nl_Product2_acc_217_nl = conv_s2s_16_18(~ (input_1_rsci_idat[63:48])) +
      ({(input_1_rsci_idat[63:48]) , 2'b01});
  assign Product2_acc_217_nl = nl_Product2_acc_217_nl[17:0];
  assign Product2_acc_217_itm_17_2_1 = readslicef_18_16_2(Product2_acc_217_nl);
  assign nl_Product2_acc_1080_nl = conv_s2u_13_17(input_1_rsci_idat[95:83]) + conv_s2u_16_17(input_1_rsci_idat[95:80]);
  assign Product2_acc_1080_nl = nl_Product2_acc_1080_nl[16:0];
  assign Product2_acc_1080_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1080_nl);
  assign nl_Product2_acc_691_nl = conv_s2s_16_20(~ (input_1_rsci_idat[159:144]))
      + ({(input_1_rsci_idat[159:144]) , 4'b0001});
  assign Product2_acc_691_nl = nl_Product2_acc_691_nl[19:0];
  assign Product2_acc_691_itm_19_4_1 = readslicef_20_16_4(Product2_acc_691_nl);
  assign nl_Product2_acc_952_nl = conv_s2s_16_20(~ (input_1_rsci_idat[223:208]))
      + ({(input_1_rsci_idat[223:208]) , 4'b0001});
  assign Product2_acc_952_nl = nl_Product2_acc_952_nl[19:0];
  assign Product2_acc_952_itm_19_4_1 = readslicef_20_16_4(Product2_acc_952_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_147_nl = ~((input_1_rsci_idat[195:192]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1
      = conv_s2s_12_13(~ (input_1_rsci_idat[207:196])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_147_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_258_nl = ~((input_1_rsci_idat[98:96]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[111:99])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_258_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Product2_acc_802_nl = conv_s2s_16_18(~ (input_1_rsci_idat[191:176]))
      + ({(input_1_rsci_idat[191:176]) , 2'b01});
  assign Product2_acc_802_nl = nl_Product2_acc_802_nl[17:0];
  assign Product2_acc_802_itm_17_2_1 = readslicef_18_16_2(Product2_acc_802_nl);
  assign nl_Product2_acc_871_nl = conv_s2s_16_18(~ (input_1_rsci_idat[207:192]))
      + ({(input_1_rsci_idat[207:192]) , 2'b01});
  assign Product2_acc_871_nl = nl_Product2_acc_871_nl[17:0];
  assign Product2_acc_871_itm_17_2_1 = readslicef_18_16_2(Product2_acc_871_nl);
  assign nl_Product2_acc_122_nl = conv_s2s_16_18(~ (input_1_rsci_idat[47:32])) +
      ({(input_1_rsci_idat[47:32]) , 2'b01});
  assign Product2_acc_122_nl = nl_Product2_acc_122_nl[17:0];
  assign Product2_acc_122_itm_17_2_1 = readslicef_18_16_2(Product2_acc_122_nl);
  assign nl_Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[111:96]);
  assign Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Product2_acc_1144_nl = conv_s2u_13_17(input_1_rsci_idat[223:211]) + conv_s2u_16_17(input_1_rsci_idat[223:208]);
  assign Product2_acc_1144_nl = nl_Product2_acc_1144_nl[16:0];
  assign Product2_acc_1144_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1144_nl);
  assign nl_Product2_acc_733_nl = conv_s2s_16_18(~ (input_1_rsci_idat[175:160]))
      + ({(input_1_rsci_idat[175:160]) , 2'b01});
  assign Product2_acc_733_nl = nl_Product2_acc_733_nl[17:0];
  assign Product2_acc_733_itm_17_2_1 = readslicef_18_16_2(Product2_acc_733_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_203_nl = ~((input_1_rsci_idat[34:32]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[47:35])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_203_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Product2_acc_216_nl = conv_s2s_16_19(~ (input_1_rsci_idat[63:48])) +
      ({(input_1_rsci_idat[63:48]) , 3'b001});
  assign Product2_acc_216_nl = nl_Product2_acc_216_nl[18:0];
  assign Product2_acc_216_itm_18_3_1 = readslicef_19_16_3(Product2_acc_216_nl);
  assign Product2_acc_1291_nl =  -conv_s2s_13_14(input_1_rsci_idat[79:67]);
  assign nl_Product2_acc_285_nl = conv_s2s_17_20({Product2_acc_1291_nl , (~ (input_1_rsci_idat[66:64]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[79:64])) , 3'b001});
  assign Product2_acc_285_nl = nl_Product2_acc_285_nl[19:0];
  assign Product2_acc_285_itm_19_4_1 = readslicef_20_16_4(Product2_acc_285_nl);
  assign nl_Product2_acc_368_cse_sva_1 = conv_s2u_12_16(input_1_rsci_idat[95:84])
      - (input_1_rsci_idat[95:80]);
  assign Product2_acc_368_cse_sva_1 = nl_Product2_acc_368_cse_sva_1[15:0];
  assign Product2_acc_1302_nl =  -conv_s2s_12_13(input_1_rsci_idat[127:116]);
  assign nl_Product2_acc_1194_nl = ({(input_1_rsci_idat[127:112]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1302_nl
      , (~ (input_1_rsci_idat[115:112]))});
  assign Product2_acc_1194_nl = nl_Product2_acc_1194_nl[17:0];
  assign nl_Product2_acc_531_nl = conv_s2s_18_20(Product2_acc_1194_nl) + ({(~ (input_1_rsci_idat[127:112]))
      , 4'b0000});
  assign Product2_acc_531_nl = nl_Product2_acc_531_nl[19:0];
  assign Product2_acc_531_itm_19_4_1 = readslicef_20_16_4(Product2_acc_531_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_338_nl = ~((input_1_rsci_idat[209:208]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[223:210])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_338_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Accum2_acc_1028_cse_1 = nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      + conv_s2s_13_14({Accum2_Accum2_conc_113_12_9 , (input_1_rsci_idat[12:4])});
  assign Accum2_acc_1028_cse_1 = nl_Accum2_acc_1028_cse_1[13:0];
  assign nl_Accum2_acc_476_cse_1 = conv_s2s_13_14(input_1_rsci_idat[191:179]) + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_476_cse_1 = nl_Accum2_acc_476_cse_1[13:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_244_nl = ~((input_1_rsci_idat[82:80]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[95:83])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_244_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Product2_acc_1175_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[79:64]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[79:64]));
  assign Product2_acc_1175_nl = nl_Product2_acc_1175_nl[18:0];
  assign nl_Product2_acc_299_nl = conv_s2s_19_20(Product2_acc_1175_nl) + ({(input_1_rsci_idat[79:64])
      , 4'b0100});
  assign Product2_acc_299_nl = nl_Product2_acc_299_nl[19:0];
  assign Product2_acc_299_itm_19_4_1 = readslicef_20_16_4(Product2_acc_299_nl);
  assign Product2_acc_1297_nl =  -conv_s2s_12_13(input_1_rsci_idat[111:100]);
  assign nl_Product2_acc_1186_nl = ({(input_1_rsci_idat[111:96]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1297_nl
      , (~ (input_1_rsci_idat[99:96]))});
  assign Product2_acc_1186_nl = nl_Product2_acc_1186_nl[17:0];
  assign nl_Product2_acc_450_nl = conv_s2s_18_20(Product2_acc_1186_nl) + ({(~ (input_1_rsci_idat[111:96]))
      , 4'b0000});
  assign Product2_acc_450_nl = nl_Product2_acc_450_nl[19:0];
  assign Product2_acc_450_itm_19_4_1 = readslicef_20_16_4(Product2_acc_450_nl);
  assign nl_Product2_acc_1117_nl = conv_s2u_13_17(input_1_rsci_idat[175:163]) + conv_s2u_16_17(input_1_rsci_idat[175:160]);
  assign Product2_acc_1117_nl = nl_Product2_acc_1117_nl[16:0];
  assign Product2_acc_1117_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1117_nl);
  assign nl_Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[223:208]);
  assign Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_182_nl = ~((input_1_rsci_idat[18:16]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[31:19])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_182_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign Product2_acc_1310_nl =  -conv_s2s_14_15(input_1_rsci_idat[191:178]);
  assign nl_Product2_acc_796_nl = conv_s2s_17_19({Product2_acc_1310_nl , (~ (input_1_rsci_idat[177:176]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[191:176])) , 2'b01});
  assign Product2_acc_796_nl = nl_Product2_acc_796_nl[18:0];
  assign Product2_acc_796_itm_18_4_1 = readslicef_19_15_4(Product2_acc_796_nl);
  assign nl_Product2_acc_370_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[95:82])
      - (input_1_rsci_idat[95:80]);
  assign Product2_acc_370_cse_sva_1 = nl_Product2_acc_370_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_42_nl = ~((input_1_rsci_idat[35:32]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1 =
      conv_s2s_12_13(~ (input_1_rsci_idat[47:36])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_42_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1[12:0];
  assign Product2_acc_1299_nl =  -conv_s2s_13_14(input_1_rsci_idat[111:99]);
  assign nl_Product2_acc_476_nl = conv_s2s_17_20({Product2_acc_1299_nl , (~ (input_1_rsci_idat[98:96]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[111:96])) , 3'b001});
  assign Product2_acc_476_nl = nl_Product2_acc_476_nl[19:0];
  assign Product2_acc_476_itm_19_4_1 = readslicef_20_16_4(Product2_acc_476_nl);
  assign nl_Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[159:144]);
  assign Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Accum2_acc_1066_cse_1 = conv_s2s_15_16(input_1_rsci_idat[95:81]) + conv_s2s_15_16(input_1_rsci_idat[111:97]);
  assign Accum2_acc_1066_cse_1 = nl_Accum2_acc_1066_cse_1[15:0];
  assign nl_Product2_acc_797_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[191:179])
      - (input_1_rsci_idat[191:176]);
  assign Product2_acc_797_cse_sva_1 = nl_Product2_acc_797_cse_sva_1[15:0];
  assign nl_Product2_acc_3_nl = conv_s2u_14_16(input_1_rsci_idat[15:2]) - (input_1_rsci_idat[15:0]);
  assign Product2_acc_3_nl = nl_Product2_acc_3_nl[15:0];
  assign Product2_acc_3_itm_15_1_1 = readslicef_16_15_1(Product2_acc_3_nl);
  assign nl_Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[63:48]);
  assign Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign Product2_acc_1290_nl =  -conv_s2s_14_15(input_1_rsci_idat[79:66]);
  assign nl_Product2_acc_283_nl = conv_s2s_17_19({Product2_acc_1290_nl , (~ (input_1_rsci_idat[65:64]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[79:64])) , 2'b01});
  assign Product2_acc_283_nl = nl_Product2_acc_283_nl[18:0];
  assign Product2_acc_283_itm_18_3_1 = readslicef_19_16_3(Product2_acc_283_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_254_nl = ~((input_1_rsci_idat[97:96]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[111:98])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_254_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_245_nl = ~((input_1_rsci_idat[81:80]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[95:82])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_245_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_1101_nl = conv_s2u_13_17(input_1_rsci_idat[127:115]) + conv_s2u_16_17(input_1_rsci_idat[127:112]);
  assign Product2_acc_1101_nl = nl_Product2_acc_1101_nl[16:0];
  assign Product2_acc_1101_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1101_nl);
  assign nl_Product2_acc_204_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[63:51])
      - (input_1_rsci_idat[63:48]);
  assign Product2_acc_204_cse_sva_1 = nl_Product2_acc_204_cse_sva_1[15:0];
  assign nl_Product2_acc_367_nl = conv_s2s_16_20(~ (input_1_rsci_idat[95:80])) +
      ({(input_1_rsci_idat[95:80]) , 4'b0001});
  assign Product2_acc_367_nl = nl_Product2_acc_367_nl[19:0];
  assign Product2_acc_367_itm_19_4_1 = readslicef_20_16_4(Product2_acc_367_nl);
  assign Product2_acc_1298_nl =  -conv_s2s_14_15(input_1_rsci_idat[111:98]);
  assign nl_Product2_acc_458_nl = conv_s2s_17_19({Product2_acc_1298_nl , (~ (input_1_rsci_idat[97:96]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[111:96])) , 2'b01});
  assign Product2_acc_458_nl = nl_Product2_acc_458_nl[18:0];
  assign Product2_acc_458_itm_18_3_1 = readslicef_19_16_3(Product2_acc_458_nl);
  assign nl_Product2_acc_1208_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[175:160]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[175:160]));
  assign Product2_acc_1208_nl = nl_Product2_acc_1208_nl[18:0];
  assign nl_Product2_acc_769_nl = conv_s2s_19_20(Product2_acc_1208_nl) + ({(input_1_rsci_idat[175:160])
      , 4'b0100});
  assign Product2_acc_769_nl = nl_Product2_acc_769_nl[19:0];
  assign Product2_acc_769_itm_19_4_1 = readslicef_20_16_4(Product2_acc_769_nl);
  assign nl_Product2_acc_943_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[223:210])
      - (input_1_rsci_idat[223:208]);
  assign Product2_acc_943_cse_sva_1 = nl_Product2_acc_943_cse_sva_1[15:0];
  assign nl_Product2_acc_730_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[175:162])
      - (input_1_rsci_idat[175:160]);
  assign Product2_acc_730_cse_sva_1 = nl_Product2_acc_730_cse_sva_1[15:0];
  assign nl_Product2_acc_667_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[159:146])
      - (input_1_rsci_idat[159:144]);
  assign Product2_acc_667_cse_sva_1 = nl_Product2_acc_667_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_262_nl = ~((input_1_rsci_idat[113:112]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[127:114])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_262_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_229_nl = ~((input_1_rsci_idat[65:64]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[79:66])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_229_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_1289_nl = conv_s2s_12_13(input_1_rsci_idat[63:52]) + 13'b0000000000001;
  assign Product2_acc_1289_nl = nl_Product2_acc_1289_nl[12:0];
  assign nl_Product2_acc_1170_nl = conv_s2s_16_17(input_1_rsci_idat[63:48]) + conv_s2s_15_17({Product2_acc_1289_nl
      , (input_1_rsci_idat[51:50])});
  assign Product2_acc_1170_nl = nl_Product2_acc_1170_nl[16:0];
  assign nl_Product2_acc_238_nl = conv_s2u_17_18(Product2_acc_1170_nl) + ({(~ (input_1_rsci_idat[63:48]))
      , 2'b00});
  assign Product2_acc_238_nl = nl_Product2_acc_238_nl[17:0];
  assign Product2_acc_238_itm_17_2_1 = readslicef_18_16_2(Product2_acc_238_nl);
  assign nl_Product2_acc_455_nl = conv_s2s_16_20(~ (input_1_rsci_idat[111:96])) +
      ({(input_1_rsci_idat[111:96]) , 4'b0001});
  assign Product2_acc_455_nl = nl_Product2_acc_455_nl[19:0];
  assign Product2_acc_455_itm_19_4_1 = readslicef_20_16_4(Product2_acc_455_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_324_nl = ~((input_1_rsci_idat[194:192]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[207:195])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_324_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Product2_acc_447_nl = conv_s2u_14_16(input_1_rsci_idat[111:98]) - (input_1_rsci_idat[111:96]);
  assign Product2_acc_447_nl = nl_Product2_acc_447_nl[15:0];
  assign Product2_acc_447_itm_15_1_1 = readslicef_16_15_1(Product2_acc_447_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_162_nl = ~((input_1_rsci_idat[211:208]!=4'b0000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1
      = conv_s2s_12_13(~ (input_1_rsci_idat[223:212])) + conv_u2s_1_13(nnet_product_mult_input_t_config2_weight_t_product_nor_162_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1 = nl_nnet_product_mult_input_t_config2_weight_t_product_acc_161_cse_sva_1[12:0];
  assign Product2_acc_1283_nl =  -conv_s2s_14_15(input_1_rsci_idat[15:2]);
  assign nl_Product2_acc_nl = conv_s2s_17_19({Product2_acc_1283_nl , (~ (input_1_rsci_idat[1:0]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[15:0])) , 2'b01});
  assign Product2_acc_nl = nl_Product2_acc_nl[18:0];
  assign Product2_acc_itm_18_3_1 = readslicef_19_16_3(Product2_acc_nl);
  assign nl_Product2_acc_1286_nl = conv_s2s_12_13(input_1_rsci_idat[47:36]) + 13'b0000000000001;
  assign Product2_acc_1286_nl = nl_Product2_acc_1286_nl[12:0];
  assign nl_Product2_acc_1165_nl = conv_s2s_16_17(input_1_rsci_idat[47:32]) + conv_s2s_15_17({Product2_acc_1286_nl
      , (input_1_rsci_idat[35:34])});
  assign Product2_acc_1165_nl = nl_Product2_acc_1165_nl[16:0];
  assign nl_Product2_acc_152_nl = conv_s2u_17_18(Product2_acc_1165_nl) + ({(~ (input_1_rsci_idat[47:32]))
      , 2'b00});
  assign Product2_acc_152_nl = nl_Product2_acc_152_nl[17:0];
  assign Product2_acc_152_itm_17_2_1 = readslicef_18_16_2(Product2_acc_152_nl);
  assign nl_Product2_acc_1197_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[127:112]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[127:112]));
  assign Product2_acc_1197_nl = nl_Product2_acc_1197_nl[18:0];
  assign nl_Product2_acc_554_nl = conv_s2s_19_20(Product2_acc_1197_nl) + ({(input_1_rsci_idat[127:112])
      , 4'b0100});
  assign Product2_acc_554_nl = nl_Product2_acc_554_nl[19:0];
  assign Product2_acc_554_itm_19_4_1 = readslicef_20_16_4(Product2_acc_554_nl);
  assign nl_Product2_acc_1105_nl = conv_s2u_14_17(input_1_rsci_idat[143:130]) + conv_s2u_16_17(input_1_rsci_idat[143:128]);
  assign Product2_acc_1105_nl = nl_Product2_acc_1105_nl[16:0];
  assign Product2_acc_1105_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1105_nl);
  assign nl_Accum2_acc_399_cse_1 = conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1)
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_399_cse_1 = nl_Accum2_acc_399_cse_1[15:0];
  assign nl_Product2_acc_85_nl = conv_s2u_14_16(input_1_rsci_idat[31:18]) - (input_1_rsci_idat[31:16]);
  assign Product2_acc_85_nl = nl_Product2_acc_85_nl[15:0];
  assign Product2_acc_85_itm_15_1_1 = readslicef_16_15_1(Product2_acc_85_nl);
  assign nl_Product2_acc_1126_nl = conv_s2u_14_17(input_1_rsci_idat[191:178]) + conv_s2u_16_17(input_1_rsci_idat[191:176]);
  assign Product2_acc_1126_nl = nl_Product2_acc_1126_nl[16:0];
  assign Product2_acc_1126_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1126_nl);
  assign nl_Product2_acc_1118_nl = conv_s2u_14_17(input_1_rsci_idat[175:162]) + conv_s2u_16_17(input_1_rsci_idat[175:160]);
  assign Product2_acc_1118_nl = nl_Product2_acc_1118_nl[16:0];
  assign Product2_acc_1118_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1118_nl);
  assign nl_Product2_acc_1221_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[223:208]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[223:208]));
  assign Product2_acc_1221_nl = nl_Product2_acc_1221_nl[18:0];
  assign nl_Product2_acc_954_nl = conv_s2s_19_20(Product2_acc_1221_nl) + ({(input_1_rsci_idat[223:208])
      , 4'b0100});
  assign Product2_acc_954_nl = nl_Product2_acc_954_nl[19:0];
  assign Product2_acc_954_itm_19_4_1 = readslicef_20_16_4(Product2_acc_954_nl);
  assign nl_Product2_acc_867_cse_sva_1 = conv_s2u_14_16(input_1_rsci_idat[207:194])
      - (input_1_rsci_idat[207:192]);
  assign Product2_acc_867_cse_sva_1 = nl_Product2_acc_867_cse_sva_1[15:0];
  assign nl_Product2_acc_629_nl = conv_s2s_16_18(~ (input_1_rsci_idat[143:128]))
      + ({(input_1_rsci_idat[143:128]) , 2'b01});
  assign Product2_acc_629_nl = nl_Product2_acc_629_nl[17:0];
  assign Product2_acc_629_itm_17_3_1 = readslicef_18_15_3(Product2_acc_629_nl);
  assign nl_Accum2_acc_1120_cse_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_120_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[95:84]);
  assign Accum2_acc_1120_cse_1 = nl_Accum2_acc_1120_cse_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_nl = ~((input_1_rsci_idat[2:0]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[15:3])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[31:17])) + conv_u2s_1_16(~ (input_1_rsci_idat[16]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[223:209])) + conv_u2s_1_16(~ (input_1_rsci_idat[208]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Product2_acc_1053_nl = conv_s2u_14_17(input_1_rsci_idat[63:50]) + conv_s2u_16_17(input_1_rsci_idat[63:48]);
  assign Product2_acc_1053_nl = nl_Product2_acc_1053_nl[16:0];
  assign Product2_acc_1053_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1053_nl);
  assign nl_Product2_acc_1184_nl = (~ (input_1_rsci_idat[111:96])) + conv_s2s_14_16(input_1_rsci_idat[111:98]);
  assign Product2_acc_1184_nl = nl_Product2_acc_1184_nl[15:0];
  assign nl_Product2_acc_1084_nl = conv_s2u_16_18(Product2_acc_1184_nl) + ({(input_1_rsci_idat[111:96])
      , 2'b01});
  assign Product2_acc_1084_nl = nl_Product2_acc_1084_nl[17:0];
  assign Product2_acc_1084_itm_17_2_1 = readslicef_18_16_2(Product2_acc_1084_nl);
  assign nl_Product2_acc_1205_nl = (~ (input_1_rsci_idat[175:160])) + conv_s2s_14_16(input_1_rsci_idat[175:162]);
  assign Product2_acc_1205_nl = nl_Product2_acc_1205_nl[15:0];
  assign nl_Product2_acc_1114_nl = conv_s2u_16_18(Product2_acc_1205_nl) + ({(input_1_rsci_idat[175:160])
      , 2'b01});
  assign Product2_acc_1114_nl = nl_Product2_acc_1114_nl[17:0];
  assign Product2_acc_1114_itm_17_2_1 = readslicef_18_16_2(Product2_acc_1114_nl);
  assign nl_Product2_acc_609_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[143:131])
      - (input_1_rsci_idat[143:128]);
  assign Product2_acc_609_cse_sva_1 = nl_Product2_acc_609_cse_sva_1[15:0];
  assign Product2_acc_1305_nl =  -conv_s2s_14_15(input_1_rsci_idat[159:146]);
  assign nl_Product2_acc_666_nl = conv_s2s_17_19({Product2_acc_1305_nl , (~ (input_1_rsci_idat[145:144]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[159:144])) , 2'b01});
  assign Product2_acc_666_nl = nl_Product2_acc_666_nl[18:0];
  assign Product2_acc_666_itm_18_3_1 = readslicef_19_16_3(Product2_acc_666_nl);
  assign nl_Product2_acc_1161_nl = (~ (input_1_rsci_idat[15:0])) + conv_s2s_14_16(input_1_rsci_idat[15:2]);
  assign Product2_acc_1161_nl = nl_Product2_acc_1161_nl[15:0];
  assign nl_Product2_acc_1028_nl = conv_s2u_16_18(Product2_acc_1161_nl) + ({(input_1_rsci_idat[15:0])
      , 2'b01});
  assign Product2_acc_1028_nl = nl_Product2_acc_1028_nl[17:0];
  assign Product2_acc_1028_itm_17_2_1 = readslicef_18_16_2(Product2_acc_1028_nl);
  assign nl_Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[31:16]);
  assign Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Product2_acc_772_nl = conv_s2s_16_19(~ (input_1_rsci_idat[175:160]))
      + ({(input_1_rsci_idat[175:160]) , 3'b001});
  assign Product2_acc_772_nl = nl_Product2_acc_772_nl[18:0];
  assign Product2_acc_772_itm_18_3_1 = readslicef_19_16_3(Product2_acc_772_nl);
  assign Product2_acc_1294_nl =  -conv_s2s_14_15(input_1_rsci_idat[95:82]);
  assign nl_Product2_acc_379_nl = conv_s2s_17_19({Product2_acc_1294_nl , (~ (input_1_rsci_idat[81:80]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[95:80])) , 2'b01});
  assign Product2_acc_379_nl = nl_Product2_acc_379_nl[18:0];
  assign Product2_acc_379_itm_18_3_1 = readslicef_19_16_3(Product2_acc_379_nl);
  assign nl_Product2_acc_166_nl = conv_s2s_16_19(~ (input_1_rsci_idat[47:32])) +
      ({(input_1_rsci_idat[47:32]) , 3'b001});
  assign Product2_acc_166_nl = nl_Product2_acc_166_nl[18:0];
  assign Product2_acc_166_itm_18_3_1 = readslicef_19_16_3(Product2_acc_166_nl);
  assign Product2_acc_1293_nl =  -conv_s2s_12_13(input_1_rsci_idat[79:68]);
  assign nl_Product2_acc_1178_nl = ({(input_1_rsci_idat[79:64]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1293_nl
      , (~ (input_1_rsci_idat[67:64]))});
  assign Product2_acc_1178_nl = nl_Product2_acc_1178_nl[17:0];
  assign nl_Product2_acc_330_nl = conv_s2s_18_20(Product2_acc_1178_nl) + ({(~ (input_1_rsci_idat[79:64]))
      , 4'b0000});
  assign Product2_acc_330_nl = nl_Product2_acc_330_nl[19:0];
  assign Product2_acc_330_itm_19_4_1 = readslicef_20_16_4(Product2_acc_330_nl);
  assign nl_Product2_acc_541_nl = conv_s2s_16_20(~ (input_1_rsci_idat[127:112]))
      + ({(input_1_rsci_idat[127:112]) , 4'b0001});
  assign Product2_acc_541_nl = nl_Product2_acc_541_nl[19:0];
  assign Product2_acc_541_itm_19_4_1 = readslicef_20_16_4(Product2_acc_541_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_311_nl = ~((input_1_rsci_idat[178:176]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[191:179])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_311_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_231_nl = ~((input_1_rsci_idat[66:64]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[79:67])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_231_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Accum2_acc_1027_cse_1 = conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1);
  assign Accum2_acc_1027_cse_1 = nl_Accum2_acc_1027_cse_1[13:0];
  assign nl_Product2_acc_1187_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[111:96]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[111:96]));
  assign Product2_acc_1187_nl = nl_Product2_acc_1187_nl[18:0];
  assign nl_Product2_acc_456_nl = conv_s2s_19_20(Product2_acc_1187_nl) + ({(input_1_rsci_idat[111:96])
      , 4'b0100});
  assign Product2_acc_456_nl = nl_Product2_acc_456_nl[19:0];
  assign Product2_acc_456_itm_19_4_1 = readslicef_20_16_4(Product2_acc_456_nl);
  assign Product2_acc_1311_nl =  -conv_s2s_13_14(input_1_rsci_idat[191:179]);
  assign nl_Product2_acc_809_nl = conv_s2s_17_20({Product2_acc_1311_nl , (~ (input_1_rsci_idat[178:176]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[191:176])) , 3'b001});
  assign Product2_acc_809_nl = nl_Product2_acc_809_nl[19:0];
  assign Product2_acc_809_itm_19_4_1 = readslicef_20_16_4(Product2_acc_809_nl);
  assign nl_Accum2_acc_825_cse_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[47:36]);
  assign Accum2_acc_825_cse_1 = nl_Accum2_acc_825_cse_1[12:0];
  assign nl_Product2_acc_671_nl = conv_s2s_16_19(~ (input_1_rsci_idat[159:144]))
      + ({(input_1_rsci_idat[159:144]) , 3'b001});
  assign Product2_acc_671_nl = nl_Product2_acc_671_nl[18:0];
  assign Product2_acc_671_itm_18_3_1 = readslicef_19_16_3(Product2_acc_671_nl);
  assign nl_Product2_acc_127_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[47:35])
      - (input_1_rsci_idat[47:32]);
  assign Product2_acc_127_cse_sva_1 = nl_Product2_acc_127_cse_sva_1[15:0];
  assign nl_Product2_acc_1176_nl = (~ (input_1_rsci_idat[79:64])) + conv_s2s_14_16(input_1_rsci_idat[79:66]);
  assign Product2_acc_1176_nl = nl_Product2_acc_1176_nl[15:0];
  assign nl_Product2_acc_1072_nl = conv_s2u_16_18(Product2_acc_1176_nl) + ({(input_1_rsci_idat[79:64])
      , 2'b01});
  assign Product2_acc_1072_nl = nl_Product2_acc_1072_nl[17:0];
  assign Product2_acc_1072_itm_17_2_1 = readslicef_18_16_2(Product2_acc_1072_nl);
  assign Product2_acc_1304_nl =  -conv_s2s_14_15(input_1_rsci_idat[143:130]);
  assign nl_Product2_acc_604_nl = conv_s2s_17_19({Product2_acc_1304_nl , (~ (input_1_rsci_idat[129:128]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[143:128])) , 2'b01});
  assign Product2_acc_604_nl = nl_Product2_acc_604_nl[18:0];
  assign Product2_acc_604_itm_18_3_1 = readslicef_19_16_3(Product2_acc_604_nl);
  assign nl_Accum2_acc_426_cse_1 = Product2_acc_455_itm_19_4_1 + Product2_acc_541_itm_19_4_1;
  assign Accum2_acc_426_cse_1 = nl_Accum2_acc_426_cse_1[15:0];
  assign Product2_acc_1314_nl =  -conv_s2s_13_14(input_1_rsci_idat[223:211]);
  assign nl_Product2_acc_932_nl = conv_s2s_17_20({Product2_acc_1314_nl , (~ (input_1_rsci_idat[210:208]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[223:208])) , 3'b001});
  assign Product2_acc_932_nl = nl_Product2_acc_932_nl[19:0];
  assign Product2_acc_932_itm_19_4_1 = readslicef_20_16_4(Product2_acc_932_nl);
  assign nl_Product2_acc_214_cse_sva_1 = conv_s2u_12_16(input_1_rsci_idat[63:52])
      - (input_1_rsci_idat[63:48]);
  assign Product2_acc_214_cse_sva_1 = nl_Product2_acc_214_cse_sva_1[15:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[79:65])) + conv_u2s_1_16(~ (input_1_rsci_idat[64]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_273_nl = ~((input_1_rsci_idat[129:128]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[143:130])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_273_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_429_nl = conv_s2s_16_19(~ (input_1_rsci_idat[95:80])) +
      ({(input_1_rsci_idat[95:80]) , 3'b001});
  assign Product2_acc_429_nl = nl_Product2_acc_429_nl[18:0];
  assign Product2_acc_429_itm_18_3_1 = readslicef_19_16_3(Product2_acc_429_nl);
  assign Product2_acc_1288_nl =  -conv_s2s_14_15(input_1_rsci_idat[63:50]);
  assign nl_Product2_acc_212_nl = conv_s2s_17_19({Product2_acc_1288_nl , (~ (input_1_rsci_idat[49:48]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[63:48])) , 2'b01});
  assign Product2_acc_212_nl = nl_Product2_acc_212_nl[18:0];
  assign Product2_acc_212_itm_18_3_1 = readslicef_19_16_3(Product2_acc_212_nl);
  assign nl_Product2_acc_1066_nl = conv_s2u_13_17(input_1_rsci_idat[79:67]) + conv_s2u_16_17(input_1_rsci_idat[79:64]);
  assign Product2_acc_1066_nl = nl_Product2_acc_1066_nl[16:0];
  assign Product2_acc_1066_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1066_nl);
  assign nl_Accum2_acc_727_cse_1 = conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_727_cse_1 = nl_Accum2_acc_727_cse_1[13:0];
  assign Product2_acc_1315_nl =  -conv_s2s_14_15(input_1_rsci_idat[223:210]);
  assign nl_Product2_acc_937_nl = conv_s2s_17_19({Product2_acc_1315_nl , (~ (input_1_rsci_idat[209:208]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[223:208])) , 2'b01});
  assign Product2_acc_937_nl = nl_Product2_acc_937_nl[18:0];
  assign Product2_acc_937_itm_18_3_1 = readslicef_19_16_3(Product2_acc_937_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_261_nl = ~((input_1_rsci_idat[114:112]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[127:115])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_261_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_310_nl = ~((input_1_rsci_idat[177:176]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[191:178])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_310_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_665_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[159:147])
      - (input_1_rsci_idat[159:144]);
  assign Product2_acc_665_cse_sva_1 = nl_Product2_acc_665_cse_sva_1[15:0];
  assign nl_Product2_acc_8_nl = conv_s2s_16_19(~ (input_1_rsci_idat[15:0])) + ({(input_1_rsci_idat[15:0])
      , 3'b001});
  assign Product2_acc_8_nl = nl_Product2_acc_8_nl[18:0];
  assign Product2_acc_8_itm_18_3_1 = readslicef_19_16_3(Product2_acc_8_nl);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[63:49])) + conv_u2s_1_16(~ (input_1_rsci_idat[48]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign Product2_acc_1301_nl =  -conv_s2s_13_14(input_1_rsci_idat[127:115]);
  assign nl_Product2_acc_528_nl = conv_s2s_17_20({Product2_acc_1301_nl , (~ (input_1_rsci_idat[114:112]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[127:112])) , 3'b001});
  assign Product2_acc_528_nl = nl_Product2_acc_528_nl[19:0];
  assign Product2_acc_528_itm_19_4_1 = readslicef_20_16_4(Product2_acc_528_nl);
  assign nl_Accum2_acc_992_cse_1 = conv_s2s_13_14(input_1_rsci_idat[31:19]) + conv_s2s_13_14(input_1_rsci_idat[95:83]);
  assign Accum2_acc_992_cse_1 = nl_Accum2_acc_992_cse_1[13:0];
  assign nl_Product2_acc_727_nl = conv_s2s_16_20(~ (input_1_rsci_idat[175:160]))
      + ({(input_1_rsci_idat[175:160]) , 4'b0001});
  assign Product2_acc_727_nl = nl_Product2_acc_727_nl[19:0];
  assign Product2_acc_727_itm_19_4_1 = readslicef_20_16_4(Product2_acc_727_nl);
  assign Product2_acc_1312_nl =  -conv_s2s_14_15(input_1_rsci_idat[207:194]);
  assign nl_Product2_acc_876_nl = conv_s2s_17_19({Product2_acc_1312_nl , (~ (input_1_rsci_idat[193:192]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[207:192])) , 2'b01});
  assign Product2_acc_876_nl = nl_Product2_acc_876_nl[18:0];
  assign Product2_acc_876_itm_18_3_1 = readslicef_19_16_3(Product2_acc_876_nl);
  assign Product2_acc_1285_nl =  -conv_s2s_14_15(input_1_rsci_idat[31:18]);
  assign nl_Product2_acc_72_nl = conv_s2s_17_19({Product2_acc_1285_nl , (~ (input_1_rsci_idat[17:16]))})
      + conv_s2s_18_19({(~ (input_1_rsci_idat[31:16])) , 2'b01});
  assign Product2_acc_72_nl = nl_Product2_acc_72_nl[18:0];
  assign Product2_acc_72_itm_18_3_1 = readslicef_19_16_3(Product2_acc_72_nl);
  assign nl_Product2_acc_141_nl = conv_s2s_16_20(~ (input_1_rsci_idat[47:32])) +
      ({(input_1_rsci_idat[47:32]) , 4'b0001});
  assign Product2_acc_141_nl = nl_Product2_acc_141_nl[19:0];
  assign Product2_acc_141_itm_19_4_1 = readslicef_20_16_4(Product2_acc_141_nl);
  assign nl_Product2_acc_499_nl = conv_s2s_16_19(~ (input_1_rsci_idat[111:96])) +
      ({(input_1_rsci_idat[111:96]) , 3'b001});
  assign Product2_acc_499_nl = nl_Product2_acc_499_nl[18:0];
  assign Product2_acc_499_itm_18_3_1 = readslicef_19_16_3(Product2_acc_499_nl);
  assign nl_Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[127:112]);
  assign Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Accum2_acc_766_cse_1 = Product2_acc_601_itm_19_4_1 + Product2_acc_667_cse_sva_1;
  assign Accum2_acc_766_cse_1 = nl_Accum2_acc_766_cse_1[15:0];
  assign nl_Accum2_acc_295_cse_1 = conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_146_cse_sva_1)
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_295_cse_1 = nl_Accum2_acc_295_cse_1[13:0];
  assign nl_Product2_acc_281_nl = conv_s2s_16_20(~ (input_1_rsci_idat[79:64])) +
      ({(input_1_rsci_idat[79:64]) , 4'b0001});
  assign Product2_acc_281_nl = nl_Product2_acc_281_nl[19:0];
  assign Product2_acc_281_itm_19_4_1 = readslicef_20_16_4(Product2_acc_281_nl);
  assign nl_Product2_acc_1095_nl = conv_s2u_14_17(input_1_rsci_idat[127:114]) + conv_s2u_16_17(input_1_rsci_idat[127:112]);
  assign Product2_acc_1095_nl = nl_Product2_acc_1095_nl[16:0];
  assign Product2_acc_1095_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1095_nl);
  assign nl_Product2_acc_970_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[223:211])
      - (input_1_rsci_idat[223:208]);
  assign Product2_acc_970_cse_sva_1 = nl_Product2_acc_970_cse_sva_1[15:0];
  assign nl_Accum2_acc_447_cse_1 = conv_s2s_14_15(input_1_rsci_idat[63:50]) + conv_s2s_14_15(input_1_rsci_idat[95:82]);
  assign Accum2_acc_447_cse_1 = nl_Accum2_acc_447_cse_1[14:0];
  assign nl_Product2_acc_1125_nl = conv_s2u_13_17(input_1_rsci_idat[191:179]) + conv_s2u_16_17(input_1_rsci_idat[191:176]);
  assign Product2_acc_1125_nl = nl_Product2_acc_1125_nl[16:0];
  assign Product2_acc_1125_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1125_nl);
  assign nl_Product2_acc_538_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[127:115])
      - (input_1_rsci_idat[127:112]);
  assign Product2_acc_538_cse_sva_1 = nl_Product2_acc_538_cse_sva_1[15:0];
  assign nl_Product2_acc_191_nl = conv_s2s_16_20(~ (input_1_rsci_idat[63:48])) +
      ({(input_1_rsci_idat[63:48]) , 4'b0001});
  assign Product2_acc_191_nl = nl_Product2_acc_191_nl[19:0];
  assign Product2_acc_191_itm_19_4_1 = readslicef_20_16_4(Product2_acc_191_nl);
  assign nl_Product2_acc_1295_nl = conv_s2s_12_13(input_1_rsci_idat[95:84]) + 13'b0000000000001;
  assign Product2_acc_1295_nl = nl_Product2_acc_1295_nl[12:0];
  assign nl_Product2_acc_1182_nl = conv_s2s_16_17(input_1_rsci_idat[95:80]) + conv_s2s_15_17({Product2_acc_1295_nl
      , (input_1_rsci_idat[83:82])});
  assign Product2_acc_1182_nl = nl_Product2_acc_1182_nl[16:0];
  assign nl_Product2_acc_394_nl = conv_s2u_17_18(Product2_acc_1182_nl) + ({(~ (input_1_rsci_idat[95:80]))
      , 2'b00});
  assign Product2_acc_394_nl = nl_Product2_acc_394_nl[17:0];
  assign Product2_acc_394_itm_17_2_1 = readslicef_18_16_2(Product2_acc_394_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_220_nl = ~((input_1_rsci_idat[50:48]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[63:51])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_220_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Product2_acc_1300_nl = conv_s2s_12_13(input_1_rsci_idat[111:100]) + 13'b0000000000001;
  assign Product2_acc_1300_nl = nl_Product2_acc_1300_nl[12:0];
  assign nl_Product2_acc_1191_nl = conv_s2s_16_17(input_1_rsci_idat[111:96]) + conv_s2s_15_17({Product2_acc_1300_nl
      , (input_1_rsci_idat[99:98])});
  assign Product2_acc_1191_nl = nl_Product2_acc_1191_nl[16:0];
  assign nl_Product2_acc_492_nl = conv_s2u_17_18(Product2_acc_1191_nl) + ({(~ (input_1_rsci_idat[111:96]))
      , 2'b00});
  assign Product2_acc_492_nl = nl_Product2_acc_492_nl[17:0];
  assign Product2_acc_492_itm_17_2_1 = readslicef_18_16_2(Product2_acc_492_nl);
  assign nl_Product2_acc_1316_nl = conv_s2s_12_13(input_1_rsci_idat[223:212]) + 13'b0000000000001;
  assign Product2_acc_1316_nl = nl_Product2_acc_1316_nl[12:0];
  assign nl_Product2_acc_1218_nl = conv_s2s_16_17(input_1_rsci_idat[223:208]) + conv_s2s_15_17({Product2_acc_1316_nl
      , (input_1_rsci_idat[211:210])});
  assign Product2_acc_1218_nl = nl_Product2_acc_1218_nl[16:0];
  assign nl_Product2_acc_942_nl = conv_s2u_17_18(Product2_acc_1218_nl) + ({(~ (input_1_rsci_idat[223:208]))
      , 2'b00});
  assign Product2_acc_942_nl = nl_Product2_acc_942_nl[17:0];
  assign Product2_acc_942_itm_17_2_1 = readslicef_18_16_2(Product2_acc_942_nl);
  assign nl_Product2_acc_1079_nl = conv_s2u_14_17(input_1_rsci_idat[95:82]) + conv_s2u_16_17(input_1_rsci_idat[95:80]);
  assign Product2_acc_1079_nl = nl_Product2_acc_1079_nl[16:0];
  assign Product2_acc_1079_itm_16_1_1 = readslicef_17_16_1(Product2_acc_1079_nl);
  assign nl_Product2_acc_1166_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[47:32]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[47:32]));
  assign Product2_acc_1166_nl = nl_Product2_acc_1166_nl[18:0];
  assign nl_Product2_acc_154_nl = conv_s2s_19_20(Product2_acc_1166_nl) + ({(input_1_rsci_idat[47:32])
      , 4'b0100});
  assign Product2_acc_154_nl = nl_Product2_acc_154_nl[19:0];
  assign Product2_acc_154_itm_19_4_1 = readslicef_20_16_4(Product2_acc_154_nl);
  assign nl_Product2_acc_1303_nl = conv_s2s_12_13(input_1_rsci_idat[127:116]) + 13'b0000000000001;
  assign Product2_acc_1303_nl = nl_Product2_acc_1303_nl[12:0];
  assign nl_Product2_acc_1196_nl = conv_s2s_16_17(input_1_rsci_idat[127:112]) + conv_s2s_15_17({Product2_acc_1303_nl
      , (input_1_rsci_idat[115:114])});
  assign Product2_acc_1196_nl = nl_Product2_acc_1196_nl[16:0];
  assign nl_Product2_acc_547_nl = conv_s2u_17_18(Product2_acc_1196_nl) + ({(~ (input_1_rsci_idat[127:112]))
      , 2'b00});
  assign Product2_acc_547_nl = nl_Product2_acc_547_nl[17:0];
  assign Product2_acc_547_itm_17_2_1 = readslicef_18_16_2(Product2_acc_547_nl);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[143:129])) + conv_u2s_1_16(~ (input_1_rsci_idat[128]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign Product2_acc_1313_nl =  -conv_s2s_13_14(input_1_rsci_idat[207:195]);
  assign nl_Product2_acc_901_nl = conv_s2s_17_20({Product2_acc_1313_nl , (~ (input_1_rsci_idat[194:192]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[207:192])) , 3'b001});
  assign Product2_acc_901_nl = nl_Product2_acc_901_nl[19:0];
  assign Product2_acc_901_itm_19_4_1 = readslicef_20_16_4(Product2_acc_901_nl);
  assign nl_Product2_acc_62_nl = conv_s2s_16_19(~ (input_1_rsci_idat[31:16])) + ({(input_1_rsci_idat[31:16])
      , 3'b001});
  assign Product2_acc_62_nl = nl_Product2_acc_62_nl[18:0];
  assign Product2_acc_62_itm_18_4_1 = readslicef_19_15_4(Product2_acc_62_nl);
  assign nl_Accum2_acc_532_cse_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_73_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[15:4]);
  assign Accum2_acc_532_cse_1 = nl_Accum2_acc_532_cse_1[12:0];
  assign nl_Product2_acc_601_nl = conv_s2s_16_20(~ (input_1_rsci_idat[143:128]))
      + ({(input_1_rsci_idat[143:128]) , 4'b0001});
  assign Product2_acc_601_nl = nl_Product2_acc_601_nl[19:0];
  assign Product2_acc_601_itm_19_4_1 = readslicef_20_16_4(Product2_acc_601_nl);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[207:193])) + conv_u2s_1_16(~ (input_1_rsci_idat[192]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Product2_acc_801_nl = conv_s2s_16_19(~ (input_1_rsci_idat[191:176]))
      + ({(input_1_rsci_idat[191:176]) , 3'b001});
  assign Product2_acc_801_nl = nl_Product2_acc_801_nl[18:0];
  assign Product2_acc_801_itm_18_4_1 = readslicef_19_15_4(Product2_acc_801_nl);
  assign nl_Product2_acc_936_cse_sva_1 = conv_s2u_12_16(input_1_rsci_idat[223:212])
      - (input_1_rsci_idat[223:208]);
  assign Product2_acc_936_cse_sva_1 = nl_Product2_acc_936_cse_sva_1[15:0];
  assign nl_Accum2_acc_306_cse_1 = nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1
      + conv_s2s_12_13(input_1_rsci_idat[15:4]);
  assign Accum2_acc_306_cse_1 = nl_Accum2_acc_306_cse_1[12:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_288_nl = ~((input_1_rsci_idat[146:144]!=3'b000));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_13_14(~ (input_1_rsci_idat[159:147])) + conv_u2s_1_14(nnet_product_mult_input_t_config2_weight_t_product_nor_288_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[13:0];
  assign nl_Accum2_acc_590_cse_1 = conv_s2s_15_16(Product2_acc_370_cse_sva_1[15:1])
      + conv_s2s_15_16(Product2_acc_1042_itm_16_1_1[15:1]);
  assign Accum2_acc_590_cse_1 = nl_Accum2_acc_590_cse_1[15:0];
  assign nl_Product2_acc_1308_nl = conv_s2s_12_13(input_1_rsci_idat[175:164]) + 13'b0000000000001;
  assign Product2_acc_1308_nl = nl_Product2_acc_1308_nl[12:0];
  assign nl_Product2_acc_1207_nl = conv_s2s_16_17(input_1_rsci_idat[175:160]) + conv_s2s_15_17({Product2_acc_1308_nl
      , (input_1_rsci_idat[163:162])});
  assign Product2_acc_1207_nl = nl_Product2_acc_1207_nl[16:0];
  assign nl_Product2_acc_742_nl = conv_s2u_17_18(Product2_acc_1207_nl) + ({(~ (input_1_rsci_idat[175:160]))
      , 2'b00});
  assign Product2_acc_742_nl = nl_Product2_acc_742_nl[17:0];
  assign Product2_acc_742_itm_17_2_1 = readslicef_18_16_2(Product2_acc_742_nl);
  assign nl_Accum2_acc_534_cse_1 = conv_s2s_13_14(input_1_rsci_idat[63:51]) + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_131_cse_sva_1);
  assign Accum2_acc_534_cse_1 = nl_Accum2_acc_534_cse_1[13:0];
  assign nl_Accum2_acc_343_cse_1 = conv_s2s_14_15(Product2_acc_667_cse_sva_1[15:2])
      + conv_s2s_14_15(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_343_cse_1 = nl_Accum2_acc_343_cse_1[14:0];
  assign nl_Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      =  -(input_1_rsci_idat[47:32]);
  assign Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_183_nl = ~((input_1_rsci_idat[17:16]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[31:18])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_183_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_794_cse_sva_1 = conv_s2u_12_16(input_1_rsci_idat[191:180])
      - (input_1_rsci_idat[191:176]);
  assign Product2_acc_794_cse_sva_1 = nl_Product2_acc_794_cse_sva_1[15:0];
  assign nl_Product2_acc_1292_nl = conv_s2s_12_13(input_1_rsci_idat[79:68]) + 13'b0000000000001;
  assign Product2_acc_1292_nl = nl_Product2_acc_1292_nl[12:0];
  assign nl_Product2_acc_1174_nl = conv_s2s_16_17(input_1_rsci_idat[79:64]) + conv_s2s_15_17({Product2_acc_1292_nl
      , (input_1_rsci_idat[67:66])});
  assign Product2_acc_1174_nl = nl_Product2_acc_1174_nl[16:0];
  assign nl_Product2_acc_298_nl = conv_s2u_17_18(Product2_acc_1174_nl) + ({(~ (input_1_rsci_idat[79:64]))
      , 2'b00});
  assign Product2_acc_298_nl = nl_Product2_acc_298_nl[17:0];
  assign Product2_acc_298_itm_17_2_1 = readslicef_18_16_2(Product2_acc_298_nl);
  assign nl_Product2_acc_560_nl = conv_s2s_16_19(~ (input_1_rsci_idat[127:112]))
      + ({(input_1_rsci_idat[127:112]) , 3'b001});
  assign Product2_acc_560_nl = nl_Product2_acc_560_nl[18:0];
  assign Product2_acc_560_itm_18_3_1 = readslicef_19_16_3(Product2_acc_560_nl);
  assign Product2_acc_1306_nl =  -conv_s2s_12_13(input_1_rsci_idat[159:148]);
  assign nl_Product2_acc_1203_nl = ({(input_1_rsci_idat[159:144]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1306_nl
      , (~ (input_1_rsci_idat[147:144]))});
  assign Product2_acc_1203_nl = nl_Product2_acc_1203_nl[17:0];
  assign nl_Product2_acc_670_nl = conv_s2s_18_20(Product2_acc_1203_nl) + ({(~ (input_1_rsci_idat[159:144]))
      , 4'b0000});
  assign Product2_acc_670_nl = nl_Product2_acc_670_nl[19:0];
  assign Product2_acc_670_itm_19_4_1 = readslicef_20_16_4(Product2_acc_670_nl);
  assign nl_Product2_acc_1309_nl = conv_s2s_12_13(input_1_rsci_idat[191:180]) + 13'b0000000000001;
  assign Product2_acc_1309_nl = nl_Product2_acc_1309_nl[12:0];
  assign nl_Product2_acc_1210_nl = conv_s2s_16_17(input_1_rsci_idat[191:176]) + conv_s2s_15_17({Product2_acc_1309_nl
      , (input_1_rsci_idat[179:178])});
  assign Product2_acc_1210_nl = nl_Product2_acc_1210_nl[16:0];
  assign nl_Product2_acc_795_nl = conv_s2u_17_18(Product2_acc_1210_nl) + ({(~ (input_1_rsci_idat[191:176]))
      , 2'b00});
  assign Product2_acc_795_nl = nl_Product2_acc_795_nl[17:0];
  assign Product2_acc_795_itm_17_2_1 = readslicef_18_16_2(Product2_acc_795_nl);
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[111:97])) + conv_u2s_1_16(~ (input_1_rsci_idat[96]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Product2_acc_1200_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[159:144]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[159:144]));
  assign Product2_acc_1200_nl = nl_Product2_acc_1200_nl[18:0];
  assign nl_Product2_acc_664_nl = conv_s2s_19_20(Product2_acc_1200_nl) + ({(input_1_rsci_idat[159:144])
      , 4'b0100});
  assign Product2_acc_664_nl = nl_Product2_acc_664_nl[19:0];
  assign Product2_acc_664_itm_19_4_1 = readslicef_20_16_4(Product2_acc_664_nl);
  assign nl_Product2_acc_382_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[95:83])
      - (input_1_rsci_idat[95:80]);
  assign Product2_acc_382_cse_sva_1 = nl_Product2_acc_382_cse_sva_1[15:0];
  assign nl_Accum2_acc_635_cse_1 = conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_41_cse_sva_1);
  assign Accum2_acc_635_cse_1 = nl_Accum2_acc_635_cse_1[13:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_300_nl = ~((input_1_rsci_idat[161:160]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[175:162])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_300_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign Product2_acc_1317_nl =  -conv_s2s_12_13(input_1_rsci_idat[223:212]);
  assign nl_Product2_acc_1220_nl = ({(input_1_rsci_idat[223:208]) , 2'b01}) + conv_s2s_17_18({Product2_acc_1317_nl
      , (~ (input_1_rsci_idat[211:208]))});
  assign Product2_acc_1220_nl = nl_Product2_acc_1220_nl[17:0];
  assign nl_Product2_acc_951_nl = conv_s2s_18_20(Product2_acc_1220_nl) + ({(~ (input_1_rsci_idat[223:208]))
      , 4'b0000});
  assign Product2_acc_951_nl = nl_Product2_acc_951_nl[19:0];
  assign Product2_acc_951_itm_19_4_1 = readslicef_20_16_4(Product2_acc_951_nl);
  assign nl_Product2_acc_743_cse_sva_1 = conv_s2u_13_16(input_1_rsci_idat[175:163])
      - (input_1_rsci_idat[175:160]);
  assign Product2_acc_743_cse_sva_1 = nl_Product2_acc_743_cse_sva_1[15:0];
  assign nl_Accum2_acc_457_cse_1 = conv_s2s_14_15(input_1_rsci_idat[31:18]) + conv_s2s_14_15(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_457_cse_1 = nl_Accum2_acc_457_cse_1[14:0];
  assign nl_Product2_acc_1284_nl = conv_s2s_12_13(input_1_rsci_idat[15:4]) + 13'b0000000000001;
  assign Product2_acc_1284_nl = nl_Product2_acc_1284_nl[12:0];
  assign nl_Product2_acc_1160_nl = conv_s2s_16_17(input_1_rsci_idat[15:0]) + conv_s2s_15_17({Product2_acc_1284_nl
      , (input_1_rsci_idat[3:2])});
  assign Product2_acc_1160_nl = nl_Product2_acc_1160_nl[16:0];
  assign nl_Product2_acc_11_nl = conv_s2u_17_18(Product2_acc_1160_nl) + ({(~ (input_1_rsci_idat[15:0]))
      , 2'b00});
  assign Product2_acc_11_nl = nl_Product2_acc_11_nl[17:0];
  assign Product2_acc_11_itm_17_2_1 = readslicef_18_16_2(Product2_acc_11_nl);
  assign Product2_acc_1287_nl =  -conv_s2s_13_14(input_1_rsci_idat[63:51]);
  assign nl_Product2_acc_193_nl = conv_s2s_17_20({Product2_acc_1287_nl , (~ (input_1_rsci_idat[50:48]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[63:48])) , 3'b001});
  assign Product2_acc_193_nl = nl_Product2_acc_193_nl[19:0];
  assign Product2_acc_193_itm_19_4_1 = readslicef_20_16_4(Product2_acc_193_nl);
  assign nl_Product2_acc_459_cse_sva_1 = conv_s2u_12_16(input_1_rsci_idat[111:100])
      - (input_1_rsci_idat[111:96]);
  assign Product2_acc_459_cse_sva_1 = nl_Product2_acc_459_cse_sva_1[15:0];
  assign Product2_acc_1296_nl =  -conv_s2s_13_14(input_1_rsci_idat[95:83]);
  assign nl_Product2_acc_398_nl = conv_s2s_17_20({Product2_acc_1296_nl , (~ (input_1_rsci_idat[82:80]))})
      + conv_s2s_19_20({(~ (input_1_rsci_idat[95:80])) , 3'b001});
  assign Product2_acc_398_nl = nl_Product2_acc_398_nl[19:0];
  assign Product2_acc_398_itm_19_4_1 = readslicef_20_16_4(Product2_acc_398_nl);
  assign nl_Product2_acc_603_nl = conv_s2u_14_16(input_1_rsci_idat[143:130]) - (input_1_rsci_idat[143:128]);
  assign Product2_acc_603_nl = nl_Product2_acc_603_nl[15:0];
  assign Product2_acc_603_itm_15_1_1 = readslicef_16_15_1(Product2_acc_603_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_nor_325_nl = ~((input_1_rsci_idat[193:192]!=2'b00));
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_14_15(~ (input_1_rsci_idat[207:194])) + conv_u2s_1_15(nnet_product_mult_input_t_config2_weight_t_product_nor_325_nl);
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[14:0];
  assign nl_Product2_acc_1163_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[31:16]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[31:16]));
  assign Product2_acc_1163_nl = nl_Product2_acc_1163_nl[18:0];
  assign nl_Product2_acc_73_nl = conv_s2s_19_20(Product2_acc_1163_nl) + ({(input_1_rsci_idat[31:16])
      , 4'b0100});
  assign Product2_acc_73_nl = nl_Product2_acc_73_nl[19:0];
  assign Product2_acc_73_itm_19_4_1 = readslicef_20_16_4(Product2_acc_73_nl);
  assign nl_Product2_acc_1199_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[143:128]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[143:128]));
  assign Product2_acc_1199_nl = nl_Product2_acc_1199_nl[18:0];
  assign nl_Product2_acc_606_nl = conv_s2s_19_20(Product2_acc_1199_nl) + ({(input_1_rsci_idat[143:128])
      , 4'b0100});
  assign Product2_acc_606_nl = nl_Product2_acc_606_nl[19:0];
  assign Product2_acc_606_itm_19_4_1 = readslicef_20_16_4(Product2_acc_606_nl);
  assign nl_Product2_acc_1179_nl = conv_s2s_18_19({(~ (input_1_rsci_idat[95:80]))
      , 2'b01}) + conv_s2s_16_19(~ (input_1_rsci_idat[95:80]));
  assign Product2_acc_1179_nl = nl_Product2_acc_1179_nl[18:0];
  assign nl_Product2_acc_374_nl = conv_s2s_19_20(Product2_acc_1179_nl) + ({(input_1_rsci_idat[95:80])
      , 4'b0100});
  assign Product2_acc_374_nl = nl_Product2_acc_374_nl[19:0];
  assign Product2_acc_374_itm_19_4_1 = readslicef_20_16_4(Product2_acc_374_nl);
  assign nl_Accum2_acc_387_cse_1 = conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_98_cse_sva_1)
      + conv_s2s_13_14(nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1);
  assign Accum2_acc_387_cse_1 = nl_Accum2_acc_387_cse_1[13:0];
  assign nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = conv_s2s_15_16(~ (input_1_rsci_idat[127:113])) + conv_u2s_1_16(~ (input_1_rsci_idat[112]));
  assign nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1
      = nl_nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1[15:0];
  assign nl_Accum2_acc_285_cse_1 = conv_s2s_15_16(Product2_acc_1053_itm_16_1_1[15:1])
      + conv_s2s_15_16(Product2_acc_1338_itm_17_3_1);
  assign Accum2_acc_285_cse_1 = nl_Accum2_acc_285_cse_1[15:0];
  assign nl_Accum2_acc_261_cse_1 = conv_s2s_15_16(Product2_acc_730_cse_sva_1[15:1])
      + conv_s2s_15_16(nnet_product_mult_input_t_config2_weight_t_product_slc_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_nnet_product_mult_input_t_config2_weight_t_product_acc_cse_sva_1);
  assign Accum2_acc_261_cse_1 = nl_Accum2_acc_261_cse_1[15:0];
  assign nl_Accum2_acc_215_cse_1 = Product2_acc_867_cse_sva_1 + Product2_acc_1144_itm_16_1_1;
  assign Accum2_acc_215_cse_1 = nl_Accum2_acc_215_cse_1[15:0];
  assign nl_Product2_acc_1330_nl = conv_s2s_16_18(~ (input_1_rsci_idat[159:144]))
      + ({(input_1_rsci_idat[159:144]) , 2'b01});
  assign Product2_acc_1330_nl = nl_Product2_acc_1330_nl[17:0];
  assign Product2_acc_1330_itm_17_3_1 = readslicef_18_15_3(Product2_acc_1330_nl);
  assign nl_Product2_acc_1332_nl = conv_s2s_16_18(~ (input_1_rsci_idat[31:16])) +
      ({(input_1_rsci_idat[31:16]) , 2'b01});
  assign Product2_acc_1332_nl = nl_Product2_acc_1332_nl[17:0];
  assign Product2_acc_1332_itm_17_2_1 = readslicef_18_16_2(Product2_acc_1332_nl);
  assign nl_Accum2_Accum2_conc_111_12_7 = conv_s2u_5_6(input_1_rsci_idat[191:187])
      + 6'b111111;
  assign Accum2_Accum2_conc_111_12_7 = nl_Accum2_Accum2_conc_111_12_7[5:0];
  assign nl_Accum2_Accum2_conc_113_12_9 = conv_s2u_3_4(input_1_rsci_idat[15:13])
      + 4'b1111;
  assign Accum2_Accum2_conc_113_12_9 = nl_Accum2_Accum2_conc_113_12_9[3:0];
  assign nl_Accum2_Accum2_conc_115_12_7 = conv_s2u_5_6(input_1_rsci_idat[207:203])
      + 6'b111011;
  assign Accum2_Accum2_conc_115_12_7 = nl_Accum2_Accum2_conc_115_12_7[5:0];
  assign nl_Accum2_Accum2_conc_117_12_6 = conv_s2u_6_7(input_1_rsci_idat[207:202])
      + 7'b0000011;
  assign Accum2_Accum2_conc_117_12_6 = nl_Accum2_Accum2_conc_117_12_6[6:0];
  assign nl_Accum2_Accum2_conc_119_12_6 = conv_s2u_6_7(input_1_rsci_idat[143:138])
      + 7'b1111111;
  assign Accum2_Accum2_conc_119_12_6 = nl_Accum2_Accum2_conc_119_12_6[6:0];
  assign nl_Accum2_Accum2_conc_121_12_8 = conv_s2u_4_5(input_1_rsci_idat[223:220])
      + 5'b11111;
  assign Accum2_Accum2_conc_121_12_8 = nl_Accum2_Accum2_conc_121_12_8[4:0];
  assign nl_Product2_acc_1334_nl = conv_s2s_16_18(~ (input_1_rsci_idat[127:112]))
      + ({(input_1_rsci_idat[127:112]) , 2'b01});
  assign Product2_acc_1334_nl = nl_Product2_acc_1334_nl[17:0];
  assign Product2_acc_1334_itm_17_3_1 = readslicef_18_15_3(Product2_acc_1334_nl);
  assign nl_Accum2_Accum2_conc_123_12_7 = conv_s2u_5_6(input_1_rsci_idat[159:155])
      + 6'b111101;
  assign Accum2_Accum2_conc_123_12_7 = nl_Accum2_Accum2_conc_123_12_7[5:0];
  assign nl_Accum2_Accum2_conc_125_12_6 = conv_s2u_6_7(input_1_rsci_idat[223:218])
      + 7'b1111001;
  assign Accum2_Accum2_conc_125_12_6 = nl_Accum2_Accum2_conc_125_12_6[6:0];
  assign nl_Product2_acc_1336_nl = conv_s2s_16_19(~ (input_1_rsci_idat[79:64])) +
      ({(input_1_rsci_idat[79:64]) , 3'b001});
  assign Product2_acc_1336_nl = nl_Product2_acc_1336_nl[18:0];
  assign Product2_acc_1336_itm_18_3_1 = readslicef_19_16_3(Product2_acc_1336_nl);
  assign nl_Product2_acc_1338_nl = conv_s2s_16_18(~ (input_1_rsci_idat[15:0])) +
      ({(input_1_rsci_idat[15:0]) , 2'b01});
  assign Product2_acc_1338_nl = nl_Product2_acc_1338_nl[17:0];
  assign Product2_acc_1338_itm_17_3_1 = readslicef_18_15_3(Product2_acc_1338_nl);
  assign nl_Accum2_Accum2_conc_127_12_7 = conv_s2u_5_6(input_1_rsci_idat[175:171])
      + 6'b111101;
  assign Accum2_Accum2_conc_127_12_7 = nl_Accum2_Accum2_conc_127_12_7[5:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_not_279 = ~(((nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_235_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_235_nl = nl_Product2_1_acc_235_nl[11:0];
  assign Product2_1_acc_235_itm_11_3_1 = readslicef_12_9_3(Product2_1_acc_235_nl);
  assign nl_Product2_1_acc_386_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_386_nl = nl_Product2_1_acc_386_nl[10:0];
  assign Product2_1_acc_386_itm_10_2_1 = readslicef_11_9_2(Product2_1_acc_386_nl);
  assign nl_Product2_1_acc_383_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_383_nl = nl_Product2_1_acc_383_nl[10:0];
  assign Product2_1_acc_383_itm_10_2_1 = readslicef_11_9_2(Product2_1_acc_383_nl);
  assign Product2_1_not_911 = ~(((nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_nl = ~(((Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_385_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_nl}) + 11'b00000000001;
  assign Product2_1_acc_385_nl = nl_Product2_1_acc_385_nl[10:0];
  assign Product2_1_acc_385_itm_10_2_1 = readslicef_11_9_2(Product2_1_acc_385_nl);
  assign Product2_1_not_941 = ~(((Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign Product2_1_not_943 = ~(((Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign Product2_1_not_949 = ~(((nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign Product2_1_not_963 = ~(((nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_acc_1110_nl = conv_s2u_14_17(input_1_rsci_idat[159:146]) + conv_s2u_16_17(input_1_rsci_idat[159:144]);
  assign Product2_acc_1110_nl = nl_Product2_acc_1110_nl[16:0];
  assign Product2_acc_1110_itm_16_2_1 = readslicef_17_15_2(Product2_acc_1110_nl);
  assign nl_Product2_acc_33_nl = conv_s2u_13_16(input_1_rsci_idat[15:3]) - (input_1_rsci_idat[15:0]);
  assign Product2_acc_33_nl = nl_Product2_acc_33_nl[15:0];
  assign Product2_acc_33_itm_15_1_1 = readslicef_16_15_1(Product2_acc_33_nl);
  assign nl_Accum2_Accum2_conc_129_12_8 = (nnet_product_mult_input_t_config2_weight_t_product_acc_14_cse_sva_1[12:8])
      + 5'b11111;
  assign Accum2_Accum2_conc_129_12_8 = nl_Accum2_Accum2_conc_129_12_8[4:0];
  assign nl_Product2_acc_290_nl = conv_s2u_13_16(input_1_rsci_idat[79:67]) - (input_1_rsci_idat[79:64]);
  assign Product2_acc_290_nl = nl_Product2_acc_290_nl[15:0];
  assign Product2_acc_290_itm_15_1_1 = readslicef_16_15_1(Product2_acc_290_nl);
  assign nl_Product2_acc_1147_nl = conv_s2u_14_17(input_1_rsci_idat[223:210]) + conv_s2u_16_17(input_1_rsci_idat[223:208]);
  assign Product2_acc_1147_nl = nl_Product2_acc_1147_nl[16:0];
  assign Product2_acc_1147_itm_16_2_1 = readslicef_17_15_2(Product2_acc_1147_nl);
  assign nl_Product2_acc_887_nl = conv_s2u_13_16(input_1_rsci_idat[207:195]) - (input_1_rsci_idat[207:192]);
  assign Product2_acc_887_nl = nl_Product2_acc_887_nl[15:0];
  assign Product2_acc_887_itm_15_1_1 = readslicef_16_15_1(Product2_acc_887_nl);
  assign nl_Accum2_acc_1648 = conv_s2s_15_16(Product2_acc_1334_itm_17_3_1) + conv_s2s_15_16(Product2_acc_1053_itm_16_1_1[15:1]);
  assign Accum2_acc_1648 = nl_Accum2_acc_1648[15:0];
  assign nl_Product2_acc_91_nl = conv_s2u_13_16(input_1_rsci_idat[31:19]) - (input_1_rsci_idat[31:16]);
  assign Product2_acc_91_nl = nl_Product2_acc_91_nl[15:0];
  assign Product2_acc_91_itm_15_1_1 = readslicef_16_15_1(Product2_acc_91_nl);
  assign nl_Product2_acc_448_nl = conv_s2u_13_16(input_1_rsci_idat[111:99]) - (input_1_rsci_idat[111:96]);
  assign Product2_acc_448_nl = nl_Product2_acc_448_nl[15:0];
  assign Product2_acc_448_itm_15_1_1 = readslicef_16_15_1(Product2_acc_448_nl);
  always @(posedge clk) begin
    if ( rst ) begin
      layer6_out_rsci_idat_14_0 <= 15'b000000000000000;
      layer6_out_rsci_idat_31_16 <= 16'b0000000000000000;
      layer6_out_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else begin
      layer6_out_rsci_idat_14_0 <= nl_layer6_out_rsci_idat_14_0[14:0];
      layer6_out_rsci_idat_31_16 <= nl_layer6_out_rsci_idat_31_16[15:0];
      layer6_out_rsci_idat_47_32 <= nl_layer6_out_rsci_idat_47_32[15:0];
    end
  end
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_8_nl = (Product2_1_acc_638_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_300_nl = conv_u2s_9_10(Product2_1_acc_638_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_8_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_300_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_300_nl[9:0];
  assign nl_Product2_1_acc_340_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_340_nl = nl_Product2_1_acc_340_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_242_nl = conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_300_nl)
      + conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_340_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_242_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_242_nl[10:0];
  assign nl_Product2_1_acc_639_nl = ({4'b1000 , (nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + 11'b00000000001;
  assign Product2_1_acc_639_nl = nl_Product2_1_acc_639_nl[10:0];
  assign nl_Product2_1_acc_640_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_640_nl = nl_Product2_1_acc_640_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_7_nl = (Product2_1_acc_636_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_299_nl = conv_u2s_9_10(Product2_1_acc_636_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_7_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_299_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_299_nl[9:0];
  assign nl_Product2_1_acc_637_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + 11'b00000000001;
  assign Product2_1_acc_637_nl = nl_Product2_1_acc_637_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_9_nl = (Product2_1_acc_641_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_301_nl = conv_u2s_9_10(Product2_1_acc_641_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_9_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_301_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_301_nl[9:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_10_nl = (Product2_1_acc_642_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_302_nl = conv_u2s_9_10(Product2_1_acc_642_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_10_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_302_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_302_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_270_nl = conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_242_nl)
      + conv_s2s_10_13(readslicef_11_10_1(Product2_1_acc_639_nl)) + conv_s2s_10_13(readslicef_11_10_1(Product2_1_acc_640_nl))
      + conv_s2s_10_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_299_nl)
      + conv_s2s_10_13(readslicef_11_10_1(Product2_1_acc_637_nl)) + conv_s2s_10_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_301_nl)
      + conv_s2s_10_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_302_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_270_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_270_nl[12:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_275_nl = conv_u2s_12_13({6'b110100
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + nnet_product_mult_layer4_t_config5_weight_t_product_acc_270_nl;
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_275_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_275_nl[12:0];
  assign nl_Product2_1_acc_300_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_300_nl = nl_Product2_1_acc_300_nl[10:0];
  assign nl_Product2_1_acc_627_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_not_911}) + 11'b00000000001;
  assign Product2_1_acc_627_nl = nl_Product2_1_acc_627_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_222_nl = conv_u2s_9_10(readslicef_11_9_2(Product2_1_acc_300_nl))
      + conv_s2s_9_10(readslicef_11_9_2(Product2_1_acc_627_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_222_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_222_nl[9:0];
  assign nl_Product2_1_acc_628_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_628_nl = nl_Product2_1_acc_628_nl[10:0];
  assign nl_Product2_1_acc_326_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_326_nl = nl_Product2_1_acc_326_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_221_nl = conv_s2s_9_10(readslicef_11_9_2(Product2_1_acc_628_nl))
      + conv_u2s_9_10(readslicef_11_9_2(Product2_1_acc_326_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_221_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_221_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_295_nl = conv_u2s_10_11(Product2_1_acc_644_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_644_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_295_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_295_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_296_nl = conv_u2s_10_11(Product2_1_acc_645_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_645_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_296_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_296_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_268_nl = conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_222_nl)
      + conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_221_nl)
      + conv_s2s_11_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_295_nl)
      + conv_s2s_11_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_296_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_268_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_268_nl[11:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_14_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_187_nl = conv_u2u_7_8(~
      (nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))
      + conv_u2u_7_8(~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_14_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_187_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_187_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_13_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_186_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_13_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_186_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_186_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_38_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_185_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:3])})
      + conv_u2u_7_8({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:3]))})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_38_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_185_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_185_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_37_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_184_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_37_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_184_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_184_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_11_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_183_nl = conv_u2u_7_8({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_7_8({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_11_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_183_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_183_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_10_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_182_nl = conv_u2u_7_8({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (layer4_out_0_9_1_lpi_1_dfm_1[8:3]))}) + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_10_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_182_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_182_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_9_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_181_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_9_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_181_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_181_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_36_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_180_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:3]))})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_36_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_180_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_180_nl[7:0];
  assign nl_Product2_1_acc_229_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_229_nl = nl_Product2_1_acc_229_nl[11:0];
  assign nl_Product2_1_acc_36_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_36_nl = nl_Product2_1_acc_36_nl[11:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_35_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_179_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_35_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_179_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_179_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_8_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_178_nl = conv_u2u_7_8({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_8_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_178_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_178_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_34_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_264_nl = conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_187_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_186_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_185_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_184_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_183_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_182_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_181_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_180_nl)
      + conv_u2u_8_12(readslicef_12_8_4(Product2_1_acc_229_nl)) + conv_u2u_8_12(Product2_1_acc_8_itm_11_2_1[9:2])
      + conv_u2u_8_12(readslicef_12_8_4(Product2_1_acc_36_nl)) + conv_u2u_8_12(Product2_1_acc_76_itm_11_4_1)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_179_nl)
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_178_nl)
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:1])})
      + conv_u2u_7_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_6_12(~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))
      + conv_u2u_1_12(nnet_product_mult_layer4_t_config5_weight_t_product_nor_34_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_264_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_264_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_272_nl = conv_s2s_12_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_268_nl)
      + conv_u2s_12_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_264_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_272_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_272_nl[13:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_nl = ~(layer4_out_0_0_lpi_1_dfm_1
      | (layer4_out_0_9_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_199_nl = conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_199_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_199_nl[8:0];
  assign nl_Product2_1_acc_174_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_174_nl = nl_Product2_1_acc_174_nl[11:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_50_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_198_nl = conv_u2u_8_9({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:2]))})
      + conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_50_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_198_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_198_nl[8:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_49_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_197_nl = conv_u2u_8_9({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_8_9({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_49_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_197_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_197_nl[8:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_263_nl = conv_u2u_9_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_199_nl)
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1])
      + conv_u2u_8_12(readslicef_12_8_4(Product2_1_acc_174_nl)) + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_9_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_198_nl)
      + conv_u2u_9_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_197_nl)
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:2]))});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_263_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_263_nl[11:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_5_nl = (Product2_1_acc_633_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_297_nl = conv_u2s_9_10(Product2_1_acc_633_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_5_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_297_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_297_nl[9:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_6_nl = (Product2_1_acc_634_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_298_nl = conv_u2s_9_10(Product2_1_acc_634_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_6_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_298_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_298_nl[9:0];
  assign nl_Product2_1_acc_624_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_624_nl = nl_Product2_1_acc_624_nl[10:0];
  assign nl_Product2_1_acc_625_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_625_nl = nl_Product2_1_acc_625_nl[10:0];
  assign nl_Product2_1_acc_629_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + 11'b00000000001;
  assign Product2_1_acc_629_nl = nl_Product2_1_acc_629_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_262_nl = conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_297_nl)
      + conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_298_nl)
      + conv_s2s_9_12(readslicef_11_9_2(Product2_1_acc_624_nl)) + conv_s2s_9_12(readslicef_11_9_2(Product2_1_acc_625_nl))
      + conv_s2s_9_12(Product2_1_acc_385_itm_10_2_1) + conv_s2s_9_12(readslicef_11_9_2(Product2_1_acc_629_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_262_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_262_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_271_nl = conv_u2s_12_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_263_nl)
      + conv_s2s_12_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_262_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_271_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_271_nl[13:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_278_nl = conv_s2s_14_15({1'b1
      , nnet_product_mult_layer4_t_config5_weight_t_product_acc_275_nl}) + conv_s2s_14_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_272_nl)
      + conv_s2s_14_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_271_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_278_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_278_nl[14:0];
  assign nl_Product2_1_acc_252_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_252_nl = nl_Product2_1_acc_252_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_227_nl = conv_u2u_9_10(readslicef_12_9_3(Product2_1_acc_252_nl))
      + conv_u2u_9_10(Product2_1_acc_235_itm_11_3_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_227_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_227_nl[9:0];
  assign nl_Product2_1_acc_622_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_622_nl = nl_Product2_1_acc_622_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_226_nl = conv_s2s_9_10(nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1)
      + conv_s2s_9_10(readslicef_11_9_2(Product2_1_acc_622_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_226_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_226_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_249_nl = conv_u2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_227_nl)
      + conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_226_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_249_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_249_nl[11:0];
  assign nl_Product2_1_acc_374_nl = conv_u2u_7_11(nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:2])
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_0});
  assign Product2_1_acc_374_nl = nl_Product2_1_acc_374_nl[10:0];
  assign nl_Product2_1_acc_631_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_631_nl = nl_Product2_1_acc_631_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_247_nl = conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_374_nl))
      + conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_631_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_247_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_247_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_267_nl = nnet_product_mult_layer4_t_config5_weight_t_product_acc_249_nl
      + conv_s2s_11_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_247_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_267_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_267_nl[11:0];
  assign nl_Product2_1_acc_34_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_34_nl = nl_Product2_1_acc_34_nl[11:0];
  assign nl_Product2_1_acc_623_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_623_nl = nl_Product2_1_acc_623_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_225_nl = conv_u2s_9_11(readslicef_12_9_3(Product2_1_acc_34_nl))
      + conv_s2s_9_11(readslicef_11_9_2(Product2_1_acc_623_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_225_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_225_nl[10:0];
  assign nl_Product2_1_acc_297_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_297_nl = nl_Product2_1_acc_297_nl[10:0];
  assign nl_Product2_1_acc_626_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_626_nl = nl_Product2_1_acc_626_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_223_nl = conv_u2s_9_10(readslicef_11_9_2(Product2_1_acc_297_nl))
      + conv_s2s_9_10(readslicef_11_9_2(Product2_1_acc_626_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_223_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_223_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_258_nl = nnet_product_mult_layer4_t_config5_weight_t_product_acc_225_nl
      + conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_223_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_258_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_258_nl[10:0];
  assign nl_Product2_1_acc_86_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_86_nl = nl_Product2_1_acc_86_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_206_nl = conv_u2u_8_9(Product2_1_acc_79_itm_11_4_1)
      + conv_u2u_8_9(readslicef_12_8_4(Product2_1_acc_86_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_206_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_206_nl[8:0];
  assign nl_Product2_1_acc_104_nl = conv_s2u_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_104_nl = nl_Product2_1_acc_104_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_205_nl = conv_u2s_8_9(readslicef_12_8_4(Product2_1_acc_104_nl))
      + conv_s2s_8_9(nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_205_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_205_nl[8:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_233_nl = conv_u2s_9_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_206_nl)
      + conv_s2s_9_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_205_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_233_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_233_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_48_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_196_nl = conv_u2u_8_9({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_8_9({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_48_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_196_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_196_nl[8:0];
  assign nl_Product2_1_acc_621_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_9
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + 11'b00000000001;
  assign Product2_1_acc_621_nl = nl_Product2_1_acc_621_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_228_nl = conv_u2s_9_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_196_nl)
      + conv_s2s_9_11(readslicef_11_9_2(Product2_1_acc_621_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_228_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_228_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_274_nl = conv_s2s_12_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_267_nl)
      + conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_258_nl)
      + conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_233_nl)
      + conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_228_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_274_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_274_nl[12:0];
  assign nl_Product2_1_acc_630_nl = ({3'b100 , (nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + 11'b00000000001;
  assign Product2_1_acc_630_nl = nl_Product2_1_acc_630_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_219_nl = conv_s2s_9_11(readslicef_11_9_2(Product2_1_acc_630_nl))
      + conv_u2s_9_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_8_1_lpi_1_dfm_1)});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_219_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_219_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_303_nl = conv_u2u_10_11(Product2_1_acc_643_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_643_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_303_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_303_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_256_nl = nnet_product_mult_layer4_t_config5_weight_t_product_acc_219_nl
      + nnet_product_mult_layer4_t_config5_weight_t_product_acc_303_nl;
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_256_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_256_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_51_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_168_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_51_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_168_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_168_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_52_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_0
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_167_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_52_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_167_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_167_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_17_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_191_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_168_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_167_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_17_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_191_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_191_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_53_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_166_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_53_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_166_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_166_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_21_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_165_nl = conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_21_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_165_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_165_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_16_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_190_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_166_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_165_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_16_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_190_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_190_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_6_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_176_nl = conv_u2u_6_7(nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])
      + conv_u2u_6_7(~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_6_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_176_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_176_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_5_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_175_nl = conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:3])})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:3]))})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_5_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_175_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_175_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_47_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_195_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_176_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_175_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_47_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_195_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_195_nl[7:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_174_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_7(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_174_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_174_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_30_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_173_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_30_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_173_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_173_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_45_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_194_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_174_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_173_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_45_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_194_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_194_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_28_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_172_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_28_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_172_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_172_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_3_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_171_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_3_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_171_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_171_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_44_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_193_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_172_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_171_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_44_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_193_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_193_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_2_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_170_nl = conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_2_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_170_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_170_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_1_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_169_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_1_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_169_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_169_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_18_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_0
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_192_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_170_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_169_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_18_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_192_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_192_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_20_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_164_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_20_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_164_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_164_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_23_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_163_nl = conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_23_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_163_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_163_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_15_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_189_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_164_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_163_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_15_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_189_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_189_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_24_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_162_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_24_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_162_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_162_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_39_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_188_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_162_nl)
      + conv_u2u_7_8(nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:2])
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_39_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_188_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_188_nl[7:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_254_nl = conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_191_nl)
      + conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_190_nl)
      + conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_195_nl)
      + conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_194_nl)
      + conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_193_nl)
      + conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_192_nl)
      + conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_189_nl)
      + conv_u2u_8_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_188_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_254_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_254_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_265_nl = conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_256_nl)
      + conv_u2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_254_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_265_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_265_nl[12:0];
  assign nl_Product2_1_acc_368_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_368_nl = nl_Product2_1_acc_368_nl[10:0];
  assign nl_Product2_1_acc_632_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_632_nl = nl_Product2_1_acc_632_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_246_nl = conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_368_nl))
      + conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_632_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_246_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_246_nl[10:0];
  assign nl_Product2_1_acc_635_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_635_nl = nl_Product2_1_acc_635_nl[10:0];
  assign nl_Product2_1_acc_303_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_303_nl = nl_Product2_1_acc_303_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_244_nl = conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_635_nl))
      + conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_303_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_244_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_244_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_273_nl = nnet_product_mult_layer4_t_config5_weight_t_product_acc_265_nl
      + conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_246_nl)
      + conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_244_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_273_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_273_nl[12:0];
  assign nl_layer6_out_rsci_idat_14_0  = nnet_product_mult_layer4_t_config5_weight_t_product_acc_278_nl
      + conv_s2s_13_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_274_nl)
      + conv_s2s_13_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_273_nl);
  assign nl_Product2_1_acc_39_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_39_nl = nl_Product2_1_acc_39_nl[11:0];
  assign nl_Product2_1_acc_517_nl = conv_s2s_9_10(nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1)
      + conv_u2s_9_10(readslicef_12_9_3(Product2_1_acc_39_nl));
  assign Product2_1_acc_517_nl = nl_Product2_1_acc_517_nl[9:0];
  assign nl_Product2_1_acc_307_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_307_nl = nl_Product2_1_acc_307_nl[10:0];
  assign nl_Product2_1_acc_123_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_123_nl = nl_Product2_1_acc_123_nl[11:0];
  assign nl_Product2_1_acc_515_nl = conv_u2u_9_10(readslicef_11_9_2(Product2_1_acc_307_nl))
      + conv_u2u_9_10(readslicef_12_9_3(Product2_1_acc_123_nl));
  assign Product2_1_acc_515_nl = nl_Product2_1_acc_515_nl[9:0];
  assign nl_Product2_1_acc_558_nl = conv_s2s_10_12(Product2_1_acc_517_nl) + conv_u2s_10_12(Product2_1_acc_515_nl);
  assign Product2_1_acc_558_nl = nl_Product2_1_acc_558_nl[11:0];
  assign nl_Product2_1_acc_488_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_0})
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1]);
  assign Product2_1_acc_488_nl = nl_Product2_1_acc_488_nl[11:0];
  assign nl_Product2_1_acc_655_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_488_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_655_nl = nl_Product2_1_acc_655_nl[10:0];
  assign nl_Product2_1_acc_489_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_489_nl = nl_Product2_1_acc_489_nl[11:0];
  assign nl_Product2_1_acc_742_nl = conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + conv_u2u_8_11(readslicef_12_8_4(Product2_1_acc_489_nl));
  assign Product2_1_acc_742_nl = nl_Product2_1_acc_742_nl[10:0];
  assign nl_Product2_1_acc_737_nl = Product2_1_acc_742_nl + 11'b01111000001;
  assign Product2_1_acc_737_nl = nl_Product2_1_acc_737_nl[10:0];
  assign nl_Product2_1_acc_591_nl = Product2_1_acc_558_nl + conv_s2s_11_12(Product2_1_acc_655_nl)
      + conv_s2s_11_12(Product2_1_acc_737_nl);
  assign Product2_1_acc_591_nl = nl_Product2_1_acc_591_nl[11:0];
  assign nl_Product2_1_acc_372_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_372_nl = nl_Product2_1_acc_372_nl[10:0];
  assign nl_Product2_1_acc_446_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_446_nl = nl_Product2_1_acc_446_nl[10:0];
  assign nl_Product2_1_acc_551_nl = conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_372_nl))
      + conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_446_nl));
  assign Product2_1_acc_551_nl = nl_Product2_1_acc_551_nl[10:0];
  assign nl_Product2_1_acc_449_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_449_nl = nl_Product2_1_acc_449_nl[10:0];
  assign nl_Product2_1_acc_279_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_279_nl = nl_Product2_1_acc_279_nl[10:0];
  assign nl_Product2_1_acc_548_nl = conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_449_nl))
      + conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_279_nl));
  assign Product2_1_acc_548_nl = nl_Product2_1_acc_548_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_279_nl = conv_u2s_10_11(Product2_1_acc_476_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_476_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_279_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_279_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_280_nl = conv_u2s_10_11(Product2_1_acc_477_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_477_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_280_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_280_nl[10:0];
  assign nl_Product2_1_acc_717_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2s_9_10(Product2_1_acc_478_itm_10_2_1);
  assign Product2_1_acc_717_nl = nl_Product2_1_acc_717_nl[9:0];
  assign nl_Product2_1_acc_648_nl = ({1'b1 , Product2_1_acc_717_nl}) + 11'b00000000001;
  assign Product2_1_acc_648_nl = nl_Product2_1_acc_648_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_281_nl = conv_u2s_10_11(Product2_1_acc_480_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_480_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_281_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_281_nl[10:0];
  assign nl_Product2_1_acc_481_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_481_nl = nl_Product2_1_acc_481_nl[11:0];
  assign nl_Product2_1_acc_741_nl = conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_8_11(readslicef_12_8_4(Product2_1_acc_481_nl));
  assign Product2_1_acc_741_nl = nl_Product2_1_acc_741_nl[10:0];
  assign nl_Product2_1_acc_736_nl = Product2_1_acc_741_nl + 11'b01111000001;
  assign Product2_1_acc_736_nl = nl_Product2_1_acc_736_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_282_nl = conv_u2s_10_11(Product2_1_acc_483_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_483_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_282_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_282_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_283_nl = conv_u2s_10_11(Product2_1_acc_484_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_484_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_283_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_283_nl[10:0];
  assign nl_Product2_1_acc_486_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_0})
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1]);
  assign Product2_1_acc_486_nl = nl_Product2_1_acc_486_nl[11:0];
  assign nl_Product2_1_acc_654_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_486_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_654_nl = nl_Product2_1_acc_654_nl[10:0];
  assign nl_Product2_1_acc_614_nl = conv_s2s_12_14(Product2_1_acc_591_nl) + conv_s2s_11_14(Product2_1_acc_551_nl)
      + conv_s2s_11_14(Product2_1_acc_548_nl) + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_279_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_280_nl)
      + conv_s2s_11_14(Product2_1_acc_648_nl) + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_281_nl)
      + conv_s2s_11_14(Product2_1_acc_736_nl) + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_282_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_283_nl)
      + conv_s2s_11_14(Product2_1_acc_654_nl);
  assign Product2_1_acc_614_nl = nl_Product2_1_acc_614_nl[13:0];
  assign nl_Product2_1_acc_115_nl = conv_s2s_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_115_nl = nl_Product2_1_acc_115_nl[12:0];
  assign nl_Product2_1_acc_457_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_457_nl = nl_Product2_1_acc_457_nl[10:0];
  assign nl_Product2_1_acc_538_nl = conv_u2s_10_12(readslicef_13_10_3(Product2_1_acc_115_nl))
      + conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_457_nl));
  assign Product2_1_acc_538_nl = nl_Product2_1_acc_538_nl[11:0];
  assign nl_Product2_1_acc_718_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_718_nl = nl_Product2_1_acc_718_nl[11:0];
  assign nl_Product2_1_acc_137_nl = ({Product2_1_acc_718_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_137_nl = nl_Product2_1_acc_137_nl[13:0];
  assign Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_2_nl = ~(((Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_460_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_2_nl}) + 11'b00000000001;
  assign Product2_1_acc_460_nl = nl_Product2_1_acc_460_nl[10:0];
  assign nl_Product2_1_acc_535_nl = conv_u2s_10_11(readslicef_14_10_4(Product2_1_acc_137_nl))
      + conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_460_nl));
  assign Product2_1_acc_535_nl = nl_Product2_1_acc_535_nl[10:0];
  assign nl_Product2_1_acc_588_nl = Product2_1_acc_538_nl + conv_s2s_11_12(Product2_1_acc_535_nl);
  assign Product2_1_acc_588_nl = nl_Product2_1_acc_588_nl[11:0];
  assign nl_Product2_1_acc_62_nl = conv_s2s_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_62_nl = nl_Product2_1_acc_62_nl[12:0];
  assign Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_1_nl = ~(((nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_453_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , Product2_1_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_1_nl}) + 11'b00000000001;
  assign Product2_1_acc_453_nl = nl_Product2_1_acc_453_nl[10:0];
  assign nl_Product2_1_acc_543_nl = conv_u2s_10_12(readslicef_13_10_3(Product2_1_acc_62_nl))
      + conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_453_nl));
  assign Product2_1_acc_543_nl = nl_Product2_1_acc_543_nl[11:0];
  assign nl_Product2_1_acc_102_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_102_nl = nl_Product2_1_acc_102_nl[11:0];
  assign nl_Product2_1_acc_456_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_456_nl = nl_Product2_1_acc_456_nl[10:0];
  assign nl_Product2_1_acc_540_nl = conv_u2s_10_12(readslicef_12_10_2(Product2_1_acc_102_nl))
      + conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_456_nl));
  assign Product2_1_acc_540_nl = nl_Product2_1_acc_540_nl[11:0];
  assign nl_Product2_1_acc_605_nl = conv_s2s_12_13(Product2_1_acc_588_nl) + conv_s2s_12_13(Product2_1_acc_543_nl)
      + conv_s2s_12_13(Product2_1_acc_540_nl);
  assign Product2_1_acc_605_nl = nl_Product2_1_acc_605_nl[12:0];
  assign nl_Product2_1_acc_352_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_352_nl = nl_Product2_1_acc_352_nl[10:0];
  assign nl_Product2_1_acc_465_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_465_nl = nl_Product2_1_acc_465_nl[10:0];
  assign nl_Product2_1_acc_528_nl = conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_352_nl))
      + conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_465_nl));
  assign Product2_1_acc_528_nl = nl_Product2_1_acc_528_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_19_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_Product2_1_acc_503_nl = conv_u2u_8_9(nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      + conv_u2u_8_9(Product2_1_acc_67_itm_11_4_1) + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_19_nl);
  assign Product2_1_acc_503_nl = nl_Product2_1_acc_503_nl[8:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_46_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_Product2_1_acc_502_nl = conv_u2u_8_9(Product2_1_acc_72_itm_11_3_1[8:1])
      + conv_u2u_8_9(Product2_1_acc_79_itm_11_4_1) + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_46_nl);
  assign Product2_1_acc_502_nl = nl_Product2_1_acc_502_nl[8:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_4_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_Product2_1_acc_492_nl = conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_4_nl);
  assign Product2_1_acc_492_nl = nl_Product2_1_acc_492_nl[6:0];
  assign nl_Product2_1_acc_491_nl = conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_6_7({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + 7'b0000001;
  assign Product2_1_acc_491_nl = nl_Product2_1_acc_491_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_12_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_Product2_1_acc_496_nl = conv_u2u_7_8(Product2_1_acc_492_nl) + conv_u2u_7_8(Product2_1_acc_491_nl)
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_12_nl);
  assign Product2_1_acc_496_nl = nl_Product2_1_acc_496_nl[7:0];
  assign nl_Product2_1_acc_495_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_1_8(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign Product2_1_acc_495_nl = nl_Product2_1_acc_495_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_7_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_Product2_1_acc_494_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(nnet_product_mult_layer4_t_config5_weight_t_product_nor_7_nl);
  assign Product2_1_acc_494_nl = nl_Product2_1_acc_494_nl[7:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_33_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_Product2_1_acc_560_nl = conv_u2u_9_11(Product2_1_acc_503_nl) + conv_u2u_9_11(Product2_1_acc_502_nl)
      + conv_u2u_8_11(Product2_1_acc_496_nl) + conv_u2u_8_11(Product2_1_acc_495_nl)
      + conv_u2u_8_11(Product2_1_acc_494_nl) + conv_u2u_7_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_6_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_1_11(nnet_product_mult_layer4_t_config5_weight_t_product_nor_33_nl);
  assign Product2_1_acc_560_nl = nl_Product2_1_acc_560_nl[10:0];
  assign nl_Product2_1_acc_587_nl = conv_s2s_11_13(Product2_1_acc_528_nl) + conv_u2s_11_13(Product2_1_acc_560_nl);
  assign Product2_1_acc_587_nl = nl_Product2_1_acc_587_nl[12:0];
  assign nl_Product2_1_acc_501_nl = conv_s2s_8_10(nnet_product_mult_layer4_t_config5_weight_t_product_slc_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_nnet_product_mult_layer4_t_config5_weight_t_product_acc_cse_sva_1)
      + conv_u2s_8_10({nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2s_1_10(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign Product2_1_acc_501_nl = nl_Product2_1_acc_501_nl[9:0];
  assign nl_Product2_1_acc_442_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_442_nl = nl_Product2_1_acc_442_nl[10:0];
  assign nl_Product2_1_acc_554_nl = conv_s2s_10_11(Product2_1_acc_501_nl) + conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_442_nl));
  assign Product2_1_acc_554_nl = nl_Product2_1_acc_554_nl[10:0];
  assign nl_Product2_1_acc_719_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_719_nl = nl_Product2_1_acc_719_nl[11:0];
  assign nl_Product2_1_acc_264_nl = ({Product2_1_acc_719_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_264_nl = nl_Product2_1_acc_264_nl[13:0];
  assign nl_Product2_1_acc_720_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_720_nl = nl_Product2_1_acc_720_nl[11:0];
  assign nl_Product2_1_acc_261_nl = ({Product2_1_acc_720_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_261_nl = nl_Product2_1_acc_261_nl[13:0];
  assign nl_Product2_1_acc_553_nl = conv_u2u_10_11(readslicef_14_10_4(Product2_1_acc_264_nl))
      + conv_u2u_10_11(readslicef_14_10_4(Product2_1_acc_261_nl));
  assign Product2_1_acc_553_nl = nl_Product2_1_acc_553_nl[10:0];
  assign nl_Product2_1_acc_584_nl = conv_s2s_11_12(Product2_1_acc_554_nl) + conv_u2s_11_12(Product2_1_acc_553_nl);
  assign Product2_1_acc_584_nl = nl_Product2_1_acc_584_nl[11:0];
  assign nl_Product2_1_acc_618_nl = conv_s2s_14_15(Product2_1_acc_614_nl) + conv_s2s_13_15(Product2_1_acc_605_nl)
      + conv_s2s_13_15(Product2_1_acc_587_nl) + conv_s2s_12_15(Product2_1_acc_584_nl);
  assign Product2_1_acc_618_nl = nl_Product2_1_acc_618_nl[14:0];
  assign nl_Product2_1_acc_721_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_721_nl = nl_Product2_1_acc_721_nl[11:0];
  assign nl_Product2_1_acc_175_nl = ({Product2_1_acc_721_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_175_nl = nl_Product2_1_acc_175_nl[13:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_2_nl = (Product2_1_acc_464_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_286_nl = conv_u2s_9_10(Product2_1_acc_464_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_2_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_286_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_286_nl[9:0];
  assign nl_Product2_1_acc_530_nl = conv_u2s_10_11(readslicef_14_10_4(Product2_1_acc_175_nl))
      + conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_286_nl);
  assign Product2_1_acc_530_nl = nl_Product2_1_acc_530_nl[10:0];
  assign nl_Product2_1_acc_192_nl = conv_s2u_11_14({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_0_lpi_1_dfm_1
      , 4'b0001});
  assign Product2_1_acc_192_nl = nl_Product2_1_acc_192_nl[13:0];
  assign nl_Product2_1_acc_350_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_0});
  assign Product2_1_acc_350_nl = nl_Product2_1_acc_350_nl[10:0];
  assign nl_Product2_1_acc_529_nl = conv_u2u_10_11(readslicef_14_10_4(Product2_1_acc_192_nl))
      + conv_u2u_10_11(readslicef_11_10_1(Product2_1_acc_350_nl));
  assign Product2_1_acc_529_nl = nl_Product2_1_acc_529_nl[10:0];
  assign nl_Product2_1_acc_575_nl = conv_s2s_11_13(Product2_1_acc_530_nl) + conv_u2s_11_13(Product2_1_acc_529_nl);
  assign Product2_1_acc_575_nl = nl_Product2_1_acc_575_nl[12:0];
  assign nl_Product2_1_acc_172_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_172_nl = nl_Product2_1_acc_172_nl[11:0];
  assign nl_Product2_1_acc_185_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_185_nl = nl_Product2_1_acc_185_nl[11:0];
  assign nl_Product2_1_acc_500_nl = conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_9({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_1_9(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign Product2_1_acc_500_nl = nl_Product2_1_acc_500_nl[8:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_43_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_Product2_1_acc_499_nl = conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_43_nl);
  assign Product2_1_acc_499_nl = nl_Product2_1_acc_499_nl[8:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_40_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_Product2_1_acc_498_nl = conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_9({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_1_9(nnet_product_mult_layer4_t_config5_weight_t_product_nor_40_nl);
  assign Product2_1_acc_498_nl = nl_Product2_1_acc_498_nl[8:0];
  assign nl_Product2_1_acc_497_nl = conv_u2u_8_9({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_1_9(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0);
  assign Product2_1_acc_497_nl = nl_Product2_1_acc_497_nl[8:0];
  assign nl_Product2_1_acc_187_nl = conv_s2u_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_0
      , 3'b001});
  assign Product2_1_acc_187_nl = nl_Product2_1_acc_187_nl[12:0];
  assign nl_Product2_1_acc_200_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_200_nl = nl_Product2_1_acc_200_nl[11:0];
  assign nl_Product2_1_acc_586_nl = conv_u2u_9_12(readslicef_12_9_3(Product2_1_acc_172_nl))
      + conv_u2u_9_12(readslicef_12_9_3(Product2_1_acc_185_nl)) + conv_u2u_9_12(Product2_1_acc_500_nl)
      + conv_u2u_9_12(Product2_1_acc_499_nl) + conv_u2u_9_12(Product2_1_acc_498_nl)
      + conv_u2u_9_12(Product2_1_acc_497_nl) + conv_u2u_9_12(readslicef_13_9_4(Product2_1_acc_187_nl))
      + conv_u2u_9_12(readslicef_12_9_3(Product2_1_acc_200_nl));
  assign Product2_1_acc_586_nl = nl_Product2_1_acc_586_nl[11:0];
  assign nl_Product2_1_acc_602_nl = conv_s2s_13_14(Product2_1_acc_575_nl) + conv_u2s_12_14(Product2_1_acc_586_nl);
  assign Product2_1_acc_602_nl = nl_Product2_1_acc_602_nl[13:0];
  assign nl_Product2_1_acc_7_nl = conv_s2u_11_14({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_0_lpi_1_dfm_1
      , 4'b0001});
  assign Product2_1_acc_7_nl = nl_Product2_1_acc_7_nl[13:0];
  assign nl_Product2_1_acc_276_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_276_nl = nl_Product2_1_acc_276_nl[10:0];
  assign nl_Product2_1_acc_549_nl = conv_u2u_10_11(readslicef_14_10_4(Product2_1_acc_7_nl))
      + conv_u2u_10_11(readslicef_11_10_1(Product2_1_acc_276_nl));
  assign Product2_1_acc_549_nl = nl_Product2_1_acc_549_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_nl = (Product2_1_acc_450_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_284_nl = conv_u2s_9_10(Product2_1_acc_450_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_284_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_284_nl[9:0];
  assign nl_Product2_1_acc_281_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_281_nl = nl_Product2_1_acc_281_nl[10:0];
  assign nl_Product2_1_acc_547_nl = conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_284_nl)
      + conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_281_nl));
  assign Product2_1_acc_547_nl = nl_Product2_1_acc_547_nl[10:0];
  assign nl_Product2_1_acc_582_nl = conv_u2s_11_13(Product2_1_acc_549_nl) + conv_s2s_11_13(Product2_1_acc_547_nl);
  assign Product2_1_acc_582_nl = nl_Product2_1_acc_582_nl[12:0];
  assign nl_Product2_1_acc_158_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_158_nl = nl_Product2_1_acc_158_nl[11:0];
  assign nl_Product2_1_acc_161_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_161_nl = nl_Product2_1_acc_161_nl[11:0];
  assign nl_Product2_1_acc_532_nl = conv_u2u_10_11(readslicef_12_10_2(Product2_1_acc_158_nl))
      + conv_u2u_10_11(readslicef_12_10_2(Product2_1_acc_161_nl));
  assign Product2_1_acc_532_nl = nl_Product2_1_acc_532_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_1_nl = (Product2_1_acc_462_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_285_nl = conv_u2s_9_10(Product2_1_acc_462_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_1_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_285_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_285_nl[9:0];
  assign nl_Product2_1_acc_338_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_338_nl = nl_Product2_1_acc_338_nl[10:0];
  assign nl_Product2_1_acc_531_nl = conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_285_nl)
      + conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_338_nl));
  assign Product2_1_acc_531_nl = nl_Product2_1_acc_531_nl[10:0];
  assign nl_Product2_1_acc_576_nl = conv_u2s_11_13(Product2_1_acc_532_nl) + conv_s2s_11_13(Product2_1_acc_531_nl);
  assign Product2_1_acc_576_nl = nl_Product2_1_acc_576_nl[12:0];
  assign nl_Product2_1_acc_31_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_31_nl = nl_Product2_1_acc_31_nl[11:0];
  assign nl_Product2_1_acc_43_nl = ({Product2_1_acc_722_cse_1 , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_43_nl = nl_Product2_1_acc_43_nl[13:0];
  assign nl_Product2_1_acc_289_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_289_nl = nl_Product2_1_acc_289_nl[10:0];
  assign nl_Product2_1_acc_56_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_56_nl = nl_Product2_1_acc_56_nl[11:0];
  assign nl_Product2_1_acc_581_nl = conv_u2u_10_12(readslicef_12_10_2(Product2_1_acc_31_nl))
      + conv_u2u_10_12(readslicef_14_10_4(Product2_1_acc_43_nl)) + conv_u2u_10_12(readslicef_11_10_1(Product2_1_acc_289_nl))
      + conv_u2u_10_12(readslicef_12_10_2(Product2_1_acc_56_nl));
  assign Product2_1_acc_581_nl = nl_Product2_1_acc_581_nl[11:0];
  assign nl_Product2_1_acc_452_nl = conv_u2s_8_10({nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_452_nl = nl_Product2_1_acc_452_nl[9:0];
  assign nl_Product2_1_acc_292_nl = conv_s2u_11_12({1'b1 , Product2_1_acc_452_nl})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_292_nl = nl_Product2_1_acc_292_nl[11:0];
  assign nl_Product2_1_acc_293_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_293_nl = nl_Product2_1_acc_293_nl[10:0];
  assign nl_Product2_1_acc_544_nl = conv_u2u_10_11(readslicef_12_10_2(Product2_1_acc_292_nl))
      + conv_u2u_10_11(readslicef_11_10_1(Product2_1_acc_293_nl));
  assign Product2_1_acc_544_nl = nl_Product2_1_acc_544_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_3_nl = (Product2_1_acc_454_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_287_nl = conv_u2s_9_10(Product2_1_acc_454_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_3_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_287_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_287_nl[9:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_4_nl = (Product2_1_acc_455_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_288_nl = conv_u2s_9_10(Product2_1_acc_455_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_4_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_288_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_288_nl[9:0];
  assign nl_Product2_1_acc_542_nl = conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_287_nl)
      + conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_288_nl);
  assign Product2_1_acc_542_nl = nl_Product2_1_acc_542_nl[10:0];
  assign nl_Product2_1_acc_580_nl = conv_u2s_11_12(Product2_1_acc_544_nl) + conv_s2s_11_12(Product2_1_acc_542_nl);
  assign Product2_1_acc_580_nl = nl_Product2_1_acc_580_nl[11:0];
  assign nl_Product2_1_acc_600_nl = conv_u2s_12_14(Product2_1_acc_581_nl) + conv_s2s_12_14(Product2_1_acc_580_nl);
  assign Product2_1_acc_600_nl = nl_Product2_1_acc_600_nl[13:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_nl
      = ~(((nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nl_Product2_1_acc_573_nl = conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_nand_nl})
      + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_573_nl = nl_Product2_1_acc_573_nl[11:0];
  assign nl_Product2_1_acc_238_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_238_nl = nl_Product2_1_acc_238_nl[11:0];
  assign nl_Product2_1_acc_519_nl = conv_s2s_9_11(Product2_1_acc_386_itm_10_2_1)
      + conv_u2s_9_11(readslicef_12_9_3(Product2_1_acc_238_nl));
  assign Product2_1_acc_519_nl = nl_Product2_1_acc_519_nl[10:0];
  assign nl_Product2_1_acc_440_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_440_nl = nl_Product2_1_acc_440_nl[10:0];
  assign nl_Product2_1_acc_227_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_227_nl = nl_Product2_1_acc_227_nl[11:0];
  assign nl_Product2_1_acc_518_nl = conv_s2s_9_11(readslicef_11_9_2(Product2_1_acc_440_nl))
      + conv_u2s_9_11(readslicef_12_9_3(Product2_1_acc_227_nl));
  assign Product2_1_acc_518_nl = nl_Product2_1_acc_518_nl[10:0];
  assign nl_Product2_1_acc_572_nl = conv_s2s_11_12(Product2_1_acc_519_nl) + conv_s2s_11_12(Product2_1_acc_518_nl);
  assign Product2_1_acc_572_nl = nl_Product2_1_acc_572_nl[11:0];
  assign nl_Product2_1_acc_597_nl = conv_u2s_12_14(Product2_1_acc_573_nl) + conv_s2s_12_14(Product2_1_acc_572_nl);
  assign Product2_1_acc_597_nl = nl_Product2_1_acc_597_nl[13:0];
  assign nl_Product2_1_acc_620_nl = conv_s2s_15_16(Product2_1_acc_618_nl) + conv_s2s_14_16(Product2_1_acc_602_nl)
      + conv_s2s_13_16(Product2_1_acc_582_nl) + conv_s2s_13_16(Product2_1_acc_576_nl)
      + conv_s2s_14_16(Product2_1_acc_600_nl) + conv_s2s_14_16(Product2_1_acc_597_nl);
  assign Product2_1_acc_620_nl = nl_Product2_1_acc_620_nl[15:0];
  assign nl_Product2_1_acc_258_nl = conv_s2u_11_14({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_0
      , 4'b0001});
  assign Product2_1_acc_258_nl = nl_Product2_1_acc_258_nl[13:0];
  assign nl_Product2_1_acc_723_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_723_nl = nl_Product2_1_acc_723_nl[11:0];
  assign nl_Product2_1_acc_248_nl = ({Product2_1_acc_723_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_248_nl = nl_Product2_1_acc_248_nl[13:0];
  assign nl_Product2_1_acc_724_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_724_nl = nl_Product2_1_acc_724_nl[11:0];
  assign nl_Product2_1_acc_231_nl = ({Product2_1_acc_724_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_231_nl = nl_Product2_1_acc_231_nl[13:0];
  assign nl_Product2_1_acc_725_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_725_nl = nl_Product2_1_acc_725_nl[11:0];
  assign nl_Product2_1_acc_6_nl = ({Product2_1_acc_725_nl , 2'b01}) + ({4'b1011 ,
      (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_6_nl = nl_Product2_1_acc_6_nl[13:0];
  assign nl_Product2_1_acc_121_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_121_nl = nl_Product2_1_acc_121_nl[11:0];
  assign nl_Product2_1_acc_125_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_125_nl = nl_Product2_1_acc_125_nl[11:0];
  assign nl_Product2_1_acc_726_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_726_nl = nl_Product2_1_acc_726_nl[11:0];
  assign nl_Product2_1_acc_126_nl = ({Product2_1_acc_726_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_126_nl = nl_Product2_1_acc_126_nl[13:0];
  assign nl_Product2_1_acc_135_nl = conv_s2u_11_14({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_0_lpi_1_dfm_1
      , 4'b0001});
  assign Product2_1_acc_135_nl = nl_Product2_1_acc_135_nl[13:0];
  assign nl_Product2_1_acc_94_nl = conv_s2u_11_14({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_0_lpi_1_dfm_1
      , 4'b0001});
  assign Product2_1_acc_94_nl = nl_Product2_1_acc_94_nl[13:0];
  assign nl_Product2_1_acc_100_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_100_nl = nl_Product2_1_acc_100_nl[11:0];
  assign nl_Product2_1_acc_313_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_313_nl = nl_Product2_1_acc_313_nl[10:0];
  assign nl_Product2_1_acc_111_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_111_nl = nl_Product2_1_acc_111_nl[11:0];
  assign nl_Product2_1_acc_610_nl = conv_u2u_9_14({nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_8_1_lpi_1_dfm_1)})
      + conv_u2u_10_14(readslicef_14_10_4(Product2_1_acc_258_nl)) + conv_u2u_10_14(readslicef_14_10_4(Product2_1_acc_248_nl))
      + conv_u2u_10_14(readslicef_14_10_4(Product2_1_acc_231_nl)) + conv_u2u_10_14(readslicef_14_10_4(Product2_1_acc_6_nl))
      + conv_u2u_10_14(readslicef_12_10_2(Product2_1_acc_121_nl)) + conv_u2u_10_14(readslicef_12_10_2(Product2_1_acc_125_nl))
      + conv_u2u_10_14(readslicef_14_10_4(Product2_1_acc_126_nl)) + conv_u2u_10_14(readslicef_14_10_4(Product2_1_acc_135_nl))
      + conv_u2u_10_14(readslicef_14_10_4(Product2_1_acc_94_nl)) + conv_u2u_10_14(readslicef_12_10_2(Product2_1_acc_100_nl))
      + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_313_nl)) + conv_u2u_10_14(readslicef_12_10_2(Product2_1_acc_111_nl))
      + conv_u2u_9_14({nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_9_lpi_1_dfm_1
      , Product2_1_acc_241_itm_11_4_1}) + conv_u2u_9_14({nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_14({nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_14({nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_8_1_lpi_1_dfm_1)})
      + conv_u2u_9_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_8_1_lpi_1_dfm_1)});
  assign Product2_1_acc_610_nl = nl_Product2_1_acc_610_nl[13:0];
  assign nl_Product2_1_acc_472_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_472_nl = nl_Product2_1_acc_472_nl[11:0];
  assign nl_Product2_1_acc_667_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_472_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_667_nl = nl_Product2_1_acc_667_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_292_nl = conv_u2s_10_11(Product2_1_acc_473_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_473_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_292_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_292_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_289_nl = conv_u2s_10_11(Product2_1_acc_466_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_466_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_289_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_289_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_290_nl = conv_u2s_10_11(Product2_1_acc_467_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_467_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_290_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_290_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_291_nl = conv_u2s_10_11(Product2_1_acc_468_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_468_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_291_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_291_nl[10:0];
  assign nl_Product2_1_acc_727_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2s_9_10(Product2_1_acc_469_itm_10_1_1[9:1]);
  assign Product2_1_acc_727_nl = nl_Product2_1_acc_727_nl[9:0];
  assign nl_Product2_1_acc_666_nl = ({1'b1 , Product2_1_acc_727_nl}) + 11'b00000000001;
  assign Product2_1_acc_666_nl = nl_Product2_1_acc_666_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_293_nl = conv_u2s_10_11(Product2_1_acc_474_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_474_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_293_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_293_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_294_nl = conv_u2s_10_11(Product2_1_acc_475_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_475_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_294_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_294_nl[10:0];
  assign nl_Product2_1_acc_608_nl = conv_s2s_11_14(Product2_1_acc_667_nl) + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_292_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_289_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_290_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_291_nl)
      + conv_s2s_11_14(Product2_1_acc_666_nl) + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_293_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_294_nl);
  assign Product2_1_acc_608_nl = nl_Product2_1_acc_608_nl[13:0];
  assign nl_Product2_1_acc_615_nl = conv_u2s_14_15(Product2_1_acc_610_nl) + conv_s2s_14_15(Product2_1_acc_608_nl);
  assign Product2_1_acc_615_nl = nl_Product2_1_acc_615_nl[14:0];
  assign nl_Product2_1_acc_355_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_355_nl = nl_Product2_1_acc_355_nl[10:0];
  assign nl_Product2_1_acc_213_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_213_nl = nl_Product2_1_acc_213_nl[11:0];
  assign nl_Product2_1_acc_461_nl = conv_u2s_8_10({nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_461_nl = nl_Product2_1_acc_461_nl[9:0];
  assign nl_Product2_1_acc_330_nl = conv_s2u_11_12({1'b1 , Product2_1_acc_461_nl})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_330_nl = nl_Product2_1_acc_330_nl[11:0];
  assign nl_Product2_1_acc_151_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_151_nl = nl_Product2_1_acc_151_nl[11:0];
  assign nl_Product2_1_acc_333_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_333_nl = nl_Product2_1_acc_333_nl[10:0];
  assign nl_Product2_1_acc_335_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_335_nl = nl_Product2_1_acc_335_nl[10:0];
  assign nl_Product2_1_acc_215_nl = conv_s2u_11_14({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_0_lpi_1_dfm_1
      , 4'b0001});
  assign Product2_1_acc_215_nl = nl_Product2_1_acc_215_nl[13:0];
  assign nl_Product2_1_acc_598_nl = conv_u2u_10_13(readslicef_11_10_1(Product2_1_acc_355_nl))
      + conv_u2u_10_13(readslicef_12_10_2(Product2_1_acc_213_nl)) + conv_u2u_10_13(readslicef_12_10_2(Product2_1_acc_330_nl))
      + conv_u2u_10_13(readslicef_12_10_2(Product2_1_acc_151_nl)) + conv_u2u_10_13(readslicef_11_10_1(Product2_1_acc_333_nl))
      + conv_u2u_10_13(readslicef_11_10_1(Product2_1_acc_335_nl)) + conv_u2u_10_13(readslicef_14_10_4(Product2_1_acc_215_nl))
      + conv_u2u_10_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1)});
  assign Product2_1_acc_598_nl = nl_Product2_1_acc_598_nl[12:0];
  assign nl_Product2_1_acc_46_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_46_nl = nl_Product2_1_acc_46_nl[11:0];
  assign nl_Product2_1_acc_516_nl = conv_u2s_9_11(readslicef_12_9_3(Product2_1_acc_46_nl))
      + conv_s2s_9_11(Product2_1_acc_383_itm_10_2_1);
  assign Product2_1_acc_516_nl = nl_Product2_1_acc_516_nl[10:0];
  assign nl_Product2_1_acc_132_nl = conv_s2u_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_132_nl = nl_Product2_1_acc_132_nl[12:0];
  assign nl_Product2_1_acc_514_nl = conv_u2s_9_10(readslicef_13_9_4(Product2_1_acc_132_nl))
      + conv_s2s_9_10(Product2_1_acc_384_itm_10_1_1[9:1]);
  assign Product2_1_acc_514_nl = nl_Product2_1_acc_514_nl[9:0];
  assign nl_Product2_1_acc_171_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_171_nl = nl_Product2_1_acc_171_nl[11:0];
  assign nl_Product2_1_acc_513_nl = conv_s2s_9_11(Product2_1_acc_385_itm_10_2_1)
      + conv_u2s_9_11(readslicef_12_9_3(Product2_1_acc_171_nl));
  assign Product2_1_acc_513_nl = nl_Product2_1_acc_513_nl[10:0];
  assign nl_Product2_1_acc_441_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_441_nl = nl_Product2_1_acc_441_nl[10:0];
  assign nl_Product2_1_acc_510_nl = conv_s2s_9_11(readslicef_11_9_2(Product2_1_acc_441_nl))
      + conv_u2s_9_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_510_nl = nl_Product2_1_acc_510_nl[10:0];
  assign nl_Product2_1_acc_596_nl = conv_s2s_11_13(Product2_1_acc_516_nl) + conv_s2s_10_13(Product2_1_acc_514_nl)
      + conv_s2s_11_13(Product2_1_acc_513_nl) + conv_s2s_11_13(Product2_1_acc_510_nl);
  assign Product2_1_acc_596_nl = nl_Product2_1_acc_596_nl[12:0];
  assign nl_Product2_1_acc_609_nl = conv_u2s_13_15(Product2_1_acc_598_nl) + conv_s2s_13_15(Product2_1_acc_596_nl);
  assign Product2_1_acc_609_nl = nl_Product2_1_acc_609_nl[14:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_27_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_Product2_1_acc_619_nl = Product2_1_acc_615_nl + Product2_1_acc_609_nl
      + ({14'b10111100000010 , nnet_product_mult_layer4_t_config5_weight_t_product_nor_27_nl});
  assign Product2_1_acc_619_nl = nl_Product2_1_acc_619_nl[14:0];
  assign nl_layer6_out_rsci_idat_31_16  = Product2_1_acc_620_nl + conv_s2s_15_16(Product2_1_acc_619_nl);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_112_nl = conv_u2u_10_12({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_112_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_112_nl[11:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_32_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_8_1_lpi_1_dfm_1[0]));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_30_nl = conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_32_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_30_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_30_nl[6:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_35_nl = conv_u2u_8_9({nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_7_9(nnet_product_mult_layer4_t_config5_weight_t_product_acc_30_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_35_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_35_nl[8:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_56_nl = conv_u2s_9_10(nnet_product_mult_layer4_t_config5_weight_t_product_acc_35_nl)
      + conv_s2s_9_10(Product2_1_acc_386_itm_10_2_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_56_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_56_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_53_nl = conv_s2s_9_10(Product2_1_acc_383_itm_10_2_1)
      + conv_u2s_9_10(Product2_1_acc_478_itm_10_2_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_53_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_53_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_111_nl = conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_56_nl)
      + conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_53_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_111_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_111_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_137_nl = conv_u2s_12_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_112_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_111_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_137_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_137_nl[13:0];
  assign nl_Product2_1_acc_21_nl = conv_s2u_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_21_nl = nl_Product2_1_acc_21_nl[12:0];
  assign nl_Product2_1_acc_164_nl = conv_s2u_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_164_nl = nl_Product2_1_acc_164_nl[12:0];
  assign nl_Product2_1_acc_168_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_168_nl = nl_Product2_1_acc_168_nl[11:0];
  assign nl_Product2_1_acc_190_nl = conv_s2u_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_190_nl = nl_Product2_1_acc_190_nl[12:0];
  assign nl_Product2_1_acc_348_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_348_nl = nl_Product2_1_acc_348_nl[10:0];
  assign nl_Product2_1_acc_218_nl = conv_s2u_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_218_nl = nl_Product2_1_acc_218_nl[12:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_144_nl = conv_u2u_9_13(readslicef_13_9_4(Product2_1_acc_21_nl))
      + conv_u2u_9_13(Product2_1_acc_72_itm_11_3_1) + conv_u2u_9_13(readslicef_13_9_4(Product2_1_acc_164_nl))
      + conv_u2u_9_13(readslicef_12_9_3(Product2_1_acc_168_nl)) + conv_u2u_9_13(readslicef_13_9_4(Product2_1_acc_190_nl))
      + conv_u2u_9_13(readslicef_11_9_2(Product2_1_acc_348_nl)) + conv_u2u_9_13(readslicef_13_9_4(Product2_1_acc_218_nl))
      + conv_u2u_9_13(nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      + conv_u2u_9_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_9_lpi_1_dfm_1
      , Product2_1_acc_241_itm_11_4_1}) + conv_u2u_9_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_13({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_8_1_lpi_1_dfm_1)})
      + conv_u2u_9_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_conc_1_pmx_8_1_lpi_1_dfm_1})
      + conv_u2u_9_13({nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_1_pmx_8_1_lpi_1_dfm_1});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_144_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_144_nl[12:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_152_nl = conv_s2s_14_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_137_nl)
      + conv_u2s_13_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_144_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_152_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_152_nl[14:0];
  assign nl_Product2_1_acc_269_nl = conv_u2u_8_11(layer4_out_0_9_1_lpi_1_dfm_1[8:1])
      + conv_u2u_10_11({layer4_out_0_9_1_lpi_1_dfm_1 , layer4_out_0_0_lpi_1_dfm_1});
  assign Product2_1_acc_269_nl = nl_Product2_1_acc_269_nl[10:0];
  assign nl_Product2_1_acc_274_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_274_nl = nl_Product2_1_acc_274_nl[10:0];
  assign nl_Product2_1_acc_18_nl = conv_s2s_11_13({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_1_pmx_0_lpi_1_dfm_1
      , 3'b001});
  assign Product2_1_acc_18_nl = nl_Product2_1_acc_18_nl[12:0];
  assign nl_Product2_1_acc_283_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_283_nl = nl_Product2_1_acc_283_nl[10:0];
  assign nl_Product2_1_acc_286_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_286_nl = nl_Product2_1_acc_286_nl[10:0];
  assign nl_Product2_1_acc_288_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_288_nl = nl_Product2_1_acc_288_nl[10:0];
  assign nl_Product2_1_acc_320_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_320_nl = nl_Product2_1_acc_320_nl[10:0];
  assign nl_Product2_1_acc_322_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_322_nl = nl_Product2_1_acc_322_nl[10:0];
  assign nl_Product2_1_acc_329_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_329_nl = nl_Product2_1_acc_329_nl[10:0];
  assign nl_Product2_1_acc_295_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_295_nl = nl_Product2_1_acc_295_nl[10:0];
  assign nl_Product2_1_acc_302_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_302_nl = nl_Product2_1_acc_302_nl[10:0];
  assign nl_Product2_1_acc_310_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_310_nl = nl_Product2_1_acc_310_nl[10:0];
  assign nl_Product2_1_acc_318_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_318_nl = nl_Product2_1_acc_318_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_151_nl = conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_269_nl))
      + conv_u2u_10_14(Product2_1_acc_469_itm_10_1_1) + conv_u2u_10_14(Product2_1_acc_8_itm_11_2_1)
      + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_274_nl)) + conv_u2u_10_14(readslicef_13_10_3(Product2_1_acc_18_nl))
      + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_283_nl)) + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_286_nl))
      + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_288_nl)) + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_320_nl))
      + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_322_nl)) + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_329_nl))
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_295_nl)) + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_302_nl))
      + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_310_nl)) + conv_u2u_10_14(readslicef_11_10_1(Product2_1_acc_318_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_151_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_151_nl[13:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_157_nl = conv_s2s_15_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_152_nl)
      + conv_u2s_14_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_151_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_157_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_157_nl[15:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_150_nl = conv_u2u_10_14({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_10_14({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_150_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_150_nl[13:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_317_nl = conv_u2s_10_11(Product2_1_acc_410_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_410_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_317_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_317_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_318_nl = conv_u2s_10_11(Product2_1_acc_411_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_411_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_318_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_318_nl[10:0];
  assign nl_Product2_1_acc_403_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_403_nl = nl_Product2_1_acc_403_nl[11:0];
  assign nl_Product2_1_acc_704_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_403_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_704_nl = nl_Product2_1_acc_704_nl[10:0];
  assign nl_Product2_1_acc_405_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_0})
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1]);
  assign Product2_1_acc_405_nl = nl_Product2_1_acc_405_nl[11:0];
  assign nl_Product2_1_acc_705_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_405_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_705_nl = nl_Product2_1_acc_705_nl[10:0];
  assign nl_Product2_1_acc_406_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_406_nl = nl_Product2_1_acc_406_nl[11:0];
  assign nl_Product2_1_acc_744_nl = conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_8_11(readslicef_12_8_4(Product2_1_acc_406_nl));
  assign Product2_1_acc_744_nl = nl_Product2_1_acc_744_nl[10:0];
  assign nl_Product2_1_acc_739_nl = Product2_1_acc_744_nl + 11'b01111000001;
  assign Product2_1_acc_739_nl = nl_Product2_1_acc_739_nl[10:0];
  assign nl_Product2_1_acc_409_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_0})
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1]);
  assign Product2_1_acc_409_nl = nl_Product2_1_acc_409_nl[11:0];
  assign nl_Product2_1_acc_708_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_409_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_708_nl = nl_Product2_1_acc_708_nl[10:0];
  assign nl_Product2_1_acc_412_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_412_nl = nl_Product2_1_acc_412_nl[11:0];
  assign nl_Product2_1_acc_745_nl = conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + conv_u2u_8_11(readslicef_12_8_4(Product2_1_acc_412_nl));
  assign Product2_1_acc_745_nl = nl_Product2_1_acc_745_nl[10:0];
  assign nl_Product2_1_acc_740_nl = Product2_1_acc_745_nl + 11'b01111000001;
  assign Product2_1_acc_740_nl = nl_Product2_1_acc_740_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_319_nl = conv_u2s_10_11(Product2_1_acc_414_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_414_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_319_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_319_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_149_nl = conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_317_nl)
      + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_318_nl)
      + conv_s2s_11_14(Product2_1_acc_704_nl) + conv_s2s_11_14(Product2_1_acc_705_nl)
      + conv_s2s_11_14(Product2_1_acc_739_nl) + conv_s2s_11_14(Product2_1_acc_708_nl)
      + conv_s2s_11_14(Product2_1_acc_740_nl) + conv_s2s_11_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_319_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_149_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_149_nl[13:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_156_nl = conv_u2s_14_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_150_nl)
      + conv_s2s_14_15(nnet_product_mult_layer4_t_config5_weight_t_product_acc_149_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_156_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_156_nl[14:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_160_nl = nnet_product_mult_layer4_t_config5_weight_t_product_acc_157_nl
      + conv_s2s_15_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_156_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_160_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_160_nl[15:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_22_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1[2:0]!=3'b000));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_312_nl = conv_u2s_10_11(Product2_1_acc_431_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_431_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_312_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_312_nl[10:0];
  assign nl_Product2_1_acc_433_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_0})
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1]);
  assign Product2_1_acc_433_nl = nl_Product2_1_acc_433_nl[11:0];
  assign nl_Product2_1_acc_696_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_433_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_696_nl = nl_Product2_1_acc_696_nl[10:0];
  assign nl_Product2_1_acc_422_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_422_nl = nl_Product2_1_acc_422_nl[11:0];
  assign nl_Product2_1_acc_687_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_422_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_687_nl = nl_Product2_1_acc_687_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_306_nl = conv_u2s_10_11(Product2_1_acc_423_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_423_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_306_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_306_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_307_nl = conv_u2s_10_11(Product2_1_acc_424_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_424_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_307_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_307_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_308_nl = conv_u2s_10_11(Product2_1_acc_425_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_425_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_308_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_308_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_304_nl = conv_u2s_10_11(Product2_1_acc_415_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_415_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_304_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_304_nl[10:0];
  assign nl_Product2_1_acc_417_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_417_nl = nl_Product2_1_acc_417_nl[11:0];
  assign nl_Product2_1_acc_683_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_417_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_683_nl = nl_Product2_1_acc_683_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_305_nl = conv_u2s_10_11(Product2_1_acc_418_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_418_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_305_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_305_nl[10:0];
  assign nl_Product2_1_acc_743_nl = conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + conv_u2u_8_11(Product2_1_acc_722_cse_1[11:4]);
  assign Product2_1_acc_743_nl = nl_Product2_1_acc_743_nl[10:0];
  assign nl_Product2_1_acc_738_nl = Product2_1_acc_743_nl + 11'b01111000001;
  assign Product2_1_acc_738_nl = nl_Product2_1_acc_738_nl[10:0];
  assign nl_Product2_1_acc_427_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_427_nl = nl_Product2_1_acc_427_nl[11:0];
  assign nl_Product2_1_acc_691_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_427_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_691_nl = nl_Product2_1_acc_691_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_309_nl = conv_u2s_10_11(Product2_1_acc_428_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_428_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_309_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_309_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_310_nl = conv_u2s_10_11(Product2_1_acc_429_itm_12_2_1[10:1])
      + ({10'b1011000000 , (Product2_1_acc_429_itm_12_2_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_310_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_310_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_311_nl = conv_u2s_10_11(Product2_1_acc_430_itm_13_3_1[10:1])
      + ({10'b1011100000 , (Product2_1_acc_430_itm_13_3_1[0])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_311_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_311_nl[10:0];
  assign nl_Product2_1_acc_435_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_0_lpi_1_dfm_1)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_0_lpi_1_dfm_1})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign Product2_1_acc_435_nl = nl_Product2_1_acc_435_nl[11:0];
  assign nl_Product2_1_acc_697_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_435_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_697_nl = nl_Product2_1_acc_697_nl[10:0];
  assign nl_Product2_1_acc_437_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_0})
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1]);
  assign Product2_1_acc_437_nl = nl_Product2_1_acc_437_nl[11:0];
  assign nl_Product2_1_acc_698_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_437_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_698_nl = nl_Product2_1_acc_698_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_159_nl = ({15'b100101101001100
      , nnet_product_mult_layer4_t_config5_weight_t_product_nor_22_nl}) + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_312_nl)
      + conv_s2s_11_16(Product2_1_acc_696_nl) + conv_s2s_11_16(Product2_1_acc_687_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_306_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_307_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_308_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_304_nl)
      + conv_s2s_11_16(Product2_1_acc_683_nl) + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_305_nl)
      + conv_s2s_11_16(Product2_1_acc_738_nl) + conv_s2s_11_16(Product2_1_acc_691_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_309_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_310_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_311_nl)
      + conv_s2s_11_16(Product2_1_acc_697_nl) + conv_s2s_11_16(Product2_1_acc_698_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_159_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_159_nl[15:0];
  assign nl_Product2_1_acc_729_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_729_nl = nl_Product2_1_acc_729_nl[11:0];
  assign nl_Product2_1_acc_177_nl = ({Product2_1_acc_729_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_177_nl = nl_Product2_1_acc_177_nl[13:0];
  assign nl_Product2_1_acc_182_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_182_nl = nl_Product2_1_acc_182_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_77_nl = conv_u2u_10_11(readslicef_14_10_4(Product2_1_acc_177_nl))
      + conv_u2u_10_11(readslicef_12_10_2(Product2_1_acc_182_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_77_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_77_nl[10:0];
  assign nl_Product2_1_acc_347_nl = conv_u2u_7_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_347_nl = nl_Product2_1_acc_347_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_11_nl = (Product2_1_acc_396_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_313_nl = conv_u2s_9_10(Product2_1_acc_396_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_11_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_313_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_313_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_76_nl = conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_347_nl))
      + conv_s2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_313_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_76_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_76_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_119_nl = conv_u2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_77_nl)
      + conv_s2s_11_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_76_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_119_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_119_nl[12:0];
  assign nl_Product2_1_acc_365_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_365_nl = nl_Product2_1_acc_365_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_128_nl = conv_u2u_8_12(Product2_1_acc_76_itm_11_4_1)
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1])
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_9_12(Product2_1_acc_235_itm_11_3_1) + conv_u2u_9_12(readslicef_11_9_2(Product2_1_acc_365_nl))
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1]))})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_8_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_128_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_128_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_145_nl = conv_s2s_13_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_119_nl)
      + conv_u2s_12_14(nnet_product_mult_layer4_t_config5_weight_t_product_acc_128_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_145_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_145_nl[13:0];
  assign nl_Product2_1_acc_387_nl = conv_u2s_8_10({nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_0_lpi_1_dfm_1)});
  assign Product2_1_acc_387_nl = nl_Product2_1_acc_387_nl[9:0];
  assign nl_Product2_1_acc_381_nl = conv_s2u_11_12({1'b1 , Product2_1_acc_387_nl})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_conc_1_pmx_0_lpi_1_dfm_1
      , 2'b01});
  assign Product2_1_acc_381_nl = nl_Product2_1_acc_381_nl[11:0];
  assign nl_Product2_1_acc_730_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_730_nl = nl_Product2_1_acc_730_nl[11:0];
  assign nl_Product2_1_acc_260_nl = ({Product2_1_acc_730_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_260_nl = nl_Product2_1_acc_260_nl[13:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_31_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_29_nl = conv_u2u_6_7({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3]))})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_31_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_29_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_29_nl[6:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_nor_29_nl = ~(nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_0_lpi_1_dfm_1
      | (nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_8_1_lpi_1_dfm_1[1:0]!=2'b00));
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_28_nl = conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_6_7({nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:3])})
      + conv_u2u_1_7(nnet_product_mult_layer4_t_config5_weight_t_product_nor_29_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_28_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_28_nl[6:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_34_nl = conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_29_nl)
      + conv_u2u_7_8(nnet_product_mult_layer4_t_config5_weight_t_product_acc_28_nl)
      + conv_u2u_1_8(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_34_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_34_nl[7:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_125_nl = conv_u2u_10_12(readslicef_12_10_2(Product2_1_acc_381_nl))
      + conv_u2u_10_12(readslicef_14_10_4(Product2_1_acc_260_nl)) + conv_u2u_9_12({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_1_pmx_8_1_lpi_1_dfm_1)})
      + conv_u2u_9_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_1_pmx_8_1_lpi_1_dfm_1)})
      + conv_u2u_9_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_1_pmx_8_1_lpi_1_dfm_1)})
      + conv_u2u_8_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_34_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_125_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_125_nl[11:0];
  assign nl_Product2_1_acc_390_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_390_nl = nl_Product2_1_acc_390_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_12_nl = (Product2_1_acc_391_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_314_nl = conv_u2s_9_10(Product2_1_acc_391_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_12_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_314_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_314_nl[9:0];
  assign nl_Product2_1_acc_392_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_392_nl = nl_Product2_1_acc_392_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_13_nl = (Product2_1_acc_393_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_315_nl = conv_u2s_9_10(Product2_1_acc_393_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_13_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_315_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_315_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_124_nl = conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_390_nl))
      + conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_314_nl)
      + conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_392_nl)) + conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_315_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_124_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_124_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_143_nl = conv_u2s_12_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_125_nl)
      + conv_s2s_12_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_124_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_143_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_143_nl[12:0];
  assign nl_Product2_1_acc_354_nl = conv_u2u_8_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_9_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_8_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_conc_1_pmx_0_lpi_1_dfm_1});
  assign Product2_1_acc_354_nl = nl_Product2_1_acc_354_nl[10:0];
  assign nl_Product2_1_acc_220_nl = conv_s2s_11_12({1'b1 , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + ({nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01});
  assign Product2_1_acc_220_nl = nl_Product2_1_acc_220_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_118_nl = conv_u2u_10_12(readslicef_11_10_1(Product2_1_acc_354_nl))
      + conv_u2u_10_12(readslicef_12_10_2(Product2_1_acc_220_nl)) + conv_u2u_10_12({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_118_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_118_nl[11:0];
  assign nl_Product2_1_acc_397_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_397_nl = nl_Product2_1_acc_397_nl[10:0];
  assign nl_Product2_1_acc_398_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_398_nl = nl_Product2_1_acc_398_nl[10:0];
  assign nnet_product_mult_layer4_t_config5_weight_t_product_and_14_nl = (Product2_1_acc_399_itm_12_2_1[1:0]==2'b11);
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_316_nl = conv_u2s_9_10(Product2_1_acc_399_itm_12_2_1[10:2])
      + ({9'b101100000 , nnet_product_mult_layer4_t_config5_weight_t_product_and_14_nl});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_316_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_316_nl[9:0];
  assign nl_Product2_1_acc_400_nl = ({3'b100 , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:1])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_400_nl = nl_Product2_1_acc_400_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_117_nl = conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_397_nl))
      + conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_398_nl)) + conv_s2s_10_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_316_nl)
      + conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_400_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_117_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_117_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_140_nl = conv_u2s_12_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_118_nl)
      + conv_s2s_12_13(nnet_product_mult_layer4_t_config5_weight_t_product_acc_117_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_140_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_140_nl[12:0];
  assign nl_Product2_1_acc_728_nl = ({nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0
      , 2'b01}) + conv_u2u_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_728_nl = nl_Product2_1_acc_728_nl[11:0];
  assign nl_Product2_1_acc_142_nl = ({Product2_1_acc_728_nl , 2'b01}) + ({4'b1011
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign Product2_1_acc_142_nl = nl_Product2_1_acc_142_nl[13:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_79_nl = conv_u2s_10_11(readslicef_14_10_4(Product2_1_acc_142_nl))
      + conv_s2s_10_11(Product2_1_acc_384_itm_10_1_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_79_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_79_nl[10:0];
  assign nl_Product2_1_acc_401_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_9)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_8_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_conc_1_pmx_lpi_1_dfm_1_0)})
      + 11'b00000000001;
  assign Product2_1_acc_401_nl = nl_Product2_1_acc_401_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_71_nl = conv_s2s_10_12(readslicef_11_10_1(Product2_1_acc_401_nl))
      + conv_u2s_10_12({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_conc_1_pmx_lpi_1_dfm_1_0)});
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_71_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_71_nl[11:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_129_nl = conv_s2s_11_12(nnet_product_mult_layer4_t_config5_weight_t_product_acc_79_nl)
      + nnet_product_mult_layer4_t_config5_weight_t_product_acc_71_nl;
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_129_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_129_nl[11:0];
  assign nl_Product2_1_acc_439_nl = ({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_9_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_0)
      , 2'b00}) + conv_u2u_10_12({nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_0})
      + conv_u2u_8_12(nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1]);
  assign Product2_1_acc_439_nl = nl_Product2_1_acc_439_nl[11:0];
  assign nl_Product2_1_acc_699_nl = ({1'b1 , (readslicef_12_10_2(Product2_1_acc_439_nl))})
      + 11'b00000000001;
  assign Product2_1_acc_699_nl = nl_Product2_1_acc_699_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_33_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_33_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_33_nl[7:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_32_nl = conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_not_279 , (~
      (nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_1_8(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_32_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_32_nl[7:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_31_nl = conv_u2u_7_8({(~
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ (nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2]))})
      + conv_u2u_7_8({nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_1_8(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_conc_1_pmx_0_lpi_1_dfm_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_31_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_31_nl[7:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_60_nl = conv_u2u_8_10(nnet_product_mult_layer4_t_config5_weight_t_product_acc_33_nl)
      + conv_u2u_8_10(nnet_product_mult_layer4_t_config5_weight_t_product_acc_32_nl)
      + conv_u2u_8_10(nnet_product_mult_layer4_t_config5_weight_t_product_acc_31_nl)
      + conv_u2u_8_10(Product2_1_acc_67_itm_11_4_1);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_60_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_60_nl[9:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_98_nl = Product2_1_acc_699_nl
      + conv_u2s_10_11(nnet_product_mult_layer4_t_config5_weight_t_product_acc_60_nl);
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_98_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_98_nl[10:0];
  assign nl_Product2_1_acc_375_nl = conv_u2u_8_11(nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1[8:1])
      + conv_u2u_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_9_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_conc_1_pmx_lpi_1_dfm_1_0});
  assign Product2_1_acc_375_nl = nl_Product2_1_acc_375_nl[10:0];
  assign nl_Product2_1_acc_389_nl = ({4'b1000 , nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1
      , (nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1[7:2])})
      + conv_u2u_10_11({(~ nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_9_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_8_1_lpi_1_dfm_1)
      , (~ nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_conc_1_pmx_0_lpi_1_dfm_1)})
      + 11'b00000000001;
  assign Product2_1_acc_389_nl = nl_Product2_1_acc_389_nl[10:0];
  assign nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_89_nl = conv_u2s_10_11(readslicef_11_10_1(Product2_1_acc_375_nl))
      + conv_s2s_10_11(readslicef_11_10_1(Product2_1_acc_389_nl));
  assign nnet_product_mult_layer4_t_config5_weight_t_product_acc_89_nl = nl_nnet_product_mult_layer4_t_config5_weight_t_product_acc_89_nl[10:0];
  assign nl_layer6_out_rsci_idat_47_32  = nnet_product_mult_layer4_t_config5_weight_t_product_acc_160_nl
      + nnet_product_mult_layer4_t_config5_weight_t_product_acc_159_nl + conv_s2s_14_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_145_nl)
      + conv_s2s_13_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_143_nl)
      + conv_s2s_13_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_140_nl)
      + conv_s2s_12_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_129_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_98_nl)
      + conv_s2s_11_16(nnet_product_mult_layer4_t_config5_weight_t_product_acc_89_nl);

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input  sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [8:0] readslicef_11_9_2;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_11_9_2 = tmp[8:0];
  end
  endfunction


  function automatic [9:0] readslicef_12_10_2;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_12_10_2 = tmp[9:0];
  end
  endfunction


  function automatic [7:0] readslicef_12_8_4;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_12_8_4 = tmp[7:0];
  end
  endfunction


  function automatic [8:0] readslicef_12_9_3;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_12_9_3 = tmp[8:0];
  end
  endfunction


  function automatic [9:0] readslicef_13_10_3;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_13_10_3 = tmp[9:0];
  end
  endfunction


  function automatic [10:0] readslicef_13_11_2;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_13_11_2 = tmp[10:0];
  end
  endfunction


  function automatic [8:0] readslicef_13_9_4;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_13_9_4 = tmp[8:0];
  end
  endfunction


  function automatic [9:0] readslicef_14_10_4;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_14_10_4 = tmp[9:0];
  end
  endfunction


  function automatic [10:0] readslicef_14_11_3;
    input [13:0] vector;
    reg [13:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_14_11_3 = tmp[10:0];
  end
  endfunction


  function automatic [14:0] readslicef_16_15_1;
    input [15:0] vector;
    reg [15:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_16_15_1 = tmp[14:0];
  end
  endfunction


  function automatic [14:0] readslicef_17_15_2;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_17_15_2 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_17_16_1;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_17_16_1 = tmp[15:0];
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [14:0] readslicef_18_15_3;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_18_15_3 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_18_16_2;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_18_16_2 = tmp[15:0];
  end
  endfunction


  function automatic [14:0] readslicef_19_15_4;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_19_15_4 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_19_16_3;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_19_16_3 = tmp[15:0];
  end
  endfunction


  function automatic [15:0] readslicef_20_16_4;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_20_16_4 = tmp[15:0];
  end
  endfunction


  function automatic [3:0] conv_s2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [4:0] conv_s2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2s_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [6:0] conv_s2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2s_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [7:0] conv_s2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_8 = {vector[6], vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_10 = {{2{vector[7]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_9_12 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_12 = {{3{vector[8]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_9_15 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_15 = {{6{vector[8]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_9_16 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_16 = {{7{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_10_12 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_12 = {{2{vector[9]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_10_13 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_13 = {{3{vector[9]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_10_14 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_14 = {{4{vector[9]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_11_13 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_13 = {{2{vector[10]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_11_14 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_14 = {{3{vector[10]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_11_16 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_16 = {{5{vector[10]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_12_14 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_14 = {{2{vector[11]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_12_15 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_15 = {{3{vector[11]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_12_16 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_16 = {{4{vector[11]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_13_15 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_15 = {{2{vector[12]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_13_16 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_16 = {{3{vector[12]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_15 = {vector[13], vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_14_16 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_16 = {{2{vector[13]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_15_16 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_16 = {vector[14], vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_15_17 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_17 = {{2{vector[14]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_16_20 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_20 = {{4{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_17_20 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_20 = {{3{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [3:0] conv_s2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2u_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2u_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2u_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_11_13 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_13 = {{2{vector[10]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_11_14 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_14 = {{3{vector[10]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2u_12_16 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_16 = {{4{vector[11]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2u_13_16 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_16 = {{3{vector[12]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_13_17 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_17 = {{4{vector[12]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2u_14_16 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_16 = {{2{vector[13]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_14_17 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_17 = {{3{vector[13]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2u_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_1_9 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_9 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_1_10 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_10 = {{9{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_1_13 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_13 = {{12{1'b0}}, vector};
  end
  endfunction


  function automatic [13:0] conv_u2s_1_14 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_14 = {{13{1'b0}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2s_1_15 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_15 = {{14{1'b0}}, vector};
  end
  endfunction


  function automatic [15:0] conv_u2s_1_16 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_16 = {{15{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_10 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_10_12 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_12 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_11_13 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_13 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2s_12_13 =  {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2s_12_14 ;
    input [11:0]  vector ;
  begin
    conv_u2s_12_14 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2s_13_15 ;
    input [12:0]  vector ;
  begin
    conv_u2s_13_15 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2s_14_15 =  {1'b0, vector};
  end
  endfunction


  function automatic [15:0] conv_u2s_14_16 ;
    input [13:0]  vector ;
  begin
    conv_u2s_14_16 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_1_7 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_7 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_1_8 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_8 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_1_9 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_9 = {{8{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_1_11 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_11 = {{10{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_1_12 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_12 = {{11{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_6_11 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_11 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_6_12 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_12 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_7_9 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_9 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_7_11 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_11 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_7_12 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_12 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_8_12 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_12 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_9_13 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_13 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_9_14 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_14 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_10_12 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_12 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_10_13 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_13 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_10_14 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_14 = {{4{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_14 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    myproject
// ------------------------------------------------------------------


module myproject (
  clk, rst, input_1_rsc_dat, layer6_out_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer6_out_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  converterBlock_myproject_core myproject_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .layer6_out_rsc_dat(layer6_out_rsc_dat)
    );
endmodule



