
//------> ./myproject_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module converterBlock_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./myproject_ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module converterBlock_ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./myproject.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
// 
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Wed Oct 26 21:54:17 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core
// ------------------------------------------------------------------


module converterBlock_myproject_core (
  clk, rst, input_1_rsc_dat, layer6_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer6_out_rsc_dat;
  input [8959:0] w2_rsc_dat;
  input [639:0] b2_rsc_dat;
  input [1919:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;


  // Interconnect Declarations
  wire [223:0] input_1_rsci_idat;
  wire [8959:0] w2_rsci_idat;
  wire [639:0] b2_rsci_idat;
  wire [1919:0] w5_rsci_idat;
  wire [14:0] b5_rsci_idat;
  reg [15:0] layer6_out_rsci_idat_47_32;
  wire [21:0] nl_layer6_out_rsci_idat_47_32;
  reg [15:0] layer6_out_rsci_idat_31_16;
  wire [21:0] nl_layer6_out_rsci_idat_31_16;
  reg [15:0] layer6_out_rsci_idat_15_0;
  wire [21:0] nl_layer6_out_rsci_idat_15_0;
  wire [15:0] Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1;
  wire [15:0] Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1;
  wire [16:0] nl_Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1;
  wire [16:0] nl_nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_0;
  wire layer4_out_conc_193_9;
  wire [7:0] layer4_out_conc_193_8_1;
  wire layer4_out_conc_193_0;
  wire layer4_out_conc_195_9;
  wire [7:0] layer4_out_conc_195_8_1;
  wire layer4_out_conc_195_0;
  wire layer4_out_conc_197_9;
  wire [7:0] layer4_out_conc_197_8_1;
  wire layer4_out_conc_197_0;
  wire layer4_out_conc_199_9;
  wire [7:0] layer4_out_conc_199_8_1;
  wire layer4_out_conc_199_0;
  wire layer4_out_conc_201_9;
  wire [7:0] layer4_out_conc_201_8_1;
  wire layer4_out_conc_201_0;
  wire layer4_out_conc_203_9;
  wire [7:0] layer4_out_conc_203_8_1;
  wire layer4_out_conc_203_0;
  wire layer4_out_conc_205_9;
  wire [7:0] layer4_out_conc_205_8_1;
  wire layer4_out_conc_205_0;
  wire layer4_out_conc_207_9;
  wire [7:0] layer4_out_conc_207_8_1;
  wire layer4_out_conc_207_0;
  wire layer4_out_conc_209_9;
  wire [7:0] layer4_out_conc_209_8_1;
  wire layer4_out_conc_209_0;
  wire layer4_out_conc_211_9;
  wire [7:0] layer4_out_conc_211_8_1;
  wire layer4_out_conc_211_0;
  wire layer4_out_conc_213_9;
  wire [7:0] layer4_out_conc_213_8_1;
  wire layer4_out_conc_213_0;
  wire layer4_out_conc_215_9;
  wire [7:0] layer4_out_conc_215_8_1;
  wire layer4_out_conc_215_0;
  wire layer4_out_conc_217_9;
  wire [7:0] layer4_out_conc_217_8_1;
  wire layer4_out_conc_217_0;
  wire layer4_out_conc_219_9;
  wire [7:0] layer4_out_conc_219_8_1;
  wire layer4_out_conc_219_0;
  wire layer4_out_conc_221_9;
  wire [7:0] layer4_out_conc_221_8_1;
  wire layer4_out_conc_221_0;
  wire layer4_out_conc_223_9;
  wire [7:0] layer4_out_conc_223_8_1;
  wire layer4_out_conc_223_0;
  wire layer4_out_conc_225_9;
  wire [7:0] layer4_out_conc_225_8_1;
  wire layer4_out_conc_225_0;
  wire layer4_out_conc_227_9;
  wire [7:0] layer4_out_conc_227_8_1;
  wire layer4_out_conc_227_0;
  wire layer4_out_conc_229_9;
  wire [7:0] layer4_out_conc_229_8_1;
  wire layer4_out_conc_229_0;
  wire layer4_out_conc_231_9;
  wire [7:0] layer4_out_conc_231_8_1;
  wire layer4_out_conc_231_0;
  wire layer4_out_conc_233_9;
  wire [7:0] layer4_out_conc_233_8_1;
  wire layer4_out_conc_233_0;
  wire layer4_out_conc_235_9;
  wire [7:0] layer4_out_conc_235_8_1;
  wire layer4_out_conc_235_0;
  wire layer4_out_conc_237_9;
  wire [7:0] layer4_out_conc_237_8_1;
  wire layer4_out_conc_237_0;
  wire layer4_out_conc_239_9;
  wire [7:0] layer4_out_conc_239_8_1;
  wire layer4_out_conc_239_0;
  wire layer4_out_conc_241_9;
  wire [7:0] layer4_out_conc_241_8_1;
  wire layer4_out_conc_241_0;
  wire layer4_out_conc_243_9;
  wire [7:0] layer4_out_conc_243_8_1;
  wire layer4_out_conc_243_0;
  wire layer4_out_conc_245_9;
  wire [7:0] layer4_out_conc_245_8_1;
  wire layer4_out_conc_245_0;
  wire layer4_out_conc_247_9;
  wire [7:0] layer4_out_conc_247_8_1;
  wire layer4_out_conc_247_0;
  wire layer4_out_conc_249_9;
  wire [7:0] layer4_out_conc_249_8_1;
  wire layer4_out_conc_249_0;
  wire layer4_out_conc_251_9;
  wire [7:0] layer4_out_conc_251_8_1;
  wire layer4_out_conc_251_0;
  wire layer4_out_conc_253_9;
  wire [7:0] layer4_out_conc_253_8_1;
  wire layer4_out_conc_253_0;
  wire layer4_out_conc_255_9;
  wire [7:0] layer4_out_conc_255_8_1;
  wire layer4_out_conc_255_0;
  wire layer4_out_conc_257_9;
  wire [7:0] layer4_out_conc_257_8_1;
  wire layer4_out_conc_257_0;
  wire layer4_out_conc_259_9;
  wire [7:0] layer4_out_conc_259_8_1;
  wire layer4_out_conc_259_0;
  wire layer4_out_conc_261_9;
  wire [7:0] layer4_out_conc_261_8_1;
  wire layer4_out_conc_261_0;
  wire layer4_out_conc_263_9;
  wire [7:0] layer4_out_conc_263_8_1;
  wire layer4_out_conc_263_0;
  wire layer4_out_conc_265_9;
  wire [7:0] layer4_out_conc_265_8_1;
  wire layer4_out_conc_265_0;
  wire layer4_out_conc_267_9;
  wire [7:0] layer4_out_conc_267_8_1;
  wire layer4_out_conc_267_0;
  wire layer4_out_conc_269_9;
  wire [7:0] layer4_out_conc_269_8_1;
  wire layer4_out_conc_269_0;
  wire layer4_out_conc_271_9;
  wire [7:0] layer4_out_conc_271_8_1;
  wire layer4_out_conc_271_0;
  wire layer4_out_conc_273_9;
  wire [7:0] layer4_out_conc_273_8_1;
  wire layer4_out_conc_273_0;
  wire layer4_out_conc_275_9;
  wire [7:0] layer4_out_conc_275_8_1;
  wire layer4_out_conc_275_0;
  wire layer4_out_conc_277_9;
  wire [7:0] layer4_out_conc_277_8_1;
  wire layer4_out_conc_277_0;
  wire layer4_out_conc_279_9;
  wire [7:0] layer4_out_conc_279_8_1;
  wire layer4_out_conc_279_0;
  wire layer4_out_conc_281_9;
  wire [7:0] layer4_out_conc_281_8_1;
  wire layer4_out_conc_281_0;
  wire layer4_out_conc_283_9;
  wire [7:0] layer4_out_conc_283_8_1;
  wire layer4_out_conc_283_0;
  wire layer4_out_conc_285_9;
  wire [7:0] layer4_out_conc_285_8_1;
  wire layer4_out_conc_285_0;
  wire layer4_out_conc_287_9;
  wire [7:0] layer4_out_conc_287_8_1;
  wire layer4_out_conc_287_0;
  wire layer4_out_conc_289_9;
  wire [7:0] layer4_out_conc_289_8_1;
  wire layer4_out_conc_289_0;
  wire layer4_out_conc_291_9;
  wire [7:0] layer4_out_conc_291_8_1;
  wire layer4_out_conc_291_0;
  wire layer4_out_conc_293_9;
  wire [7:0] layer4_out_conc_293_8_1;
  wire layer4_out_conc_293_0;
  wire layer4_out_conc_295_9;
  wire [7:0] layer4_out_conc_295_8_1;
  wire layer4_out_conc_295_0;
  wire layer4_out_conc_297_9;
  wire [7:0] layer4_out_conc_297_8_1;
  wire layer4_out_conc_297_0;
  wire layer4_out_conc_299_9;
  wire [7:0] layer4_out_conc_299_8_1;
  wire layer4_out_conc_299_0;
  wire layer4_out_conc_301_9;
  wire [7:0] layer4_out_conc_301_8_1;
  wire layer4_out_conc_301_0;
  wire layer4_out_conc_303_9;
  wire [7:0] layer4_out_conc_303_8_1;
  wire layer4_out_conc_303_0;
  wire layer4_out_conc_305_9;
  wire [7:0] layer4_out_conc_305_8_1;
  wire layer4_out_conc_305_0;
  wire layer4_out_conc_307_9;
  wire [7:0] layer4_out_conc_307_8_1;
  wire layer4_out_conc_307_0;
  wire layer4_out_conc_309_9;
  wire [7:0] layer4_out_conc_309_8_1;
  wire layer4_out_conc_309_0;
  wire layer4_out_conc_311_9;
  wire [7:0] layer4_out_conc_311_8_1;
  wire layer4_out_conc_311_0;
  wire layer4_out_conc_313_9;
  wire [7:0] layer4_out_conc_313_8_1;
  wire layer4_out_conc_313_0;
  wire layer4_out_conc_315_9;
  wire [7:0] layer4_out_conc_315_8_1;
  wire layer4_out_conc_315_0;
  wire layer4_out_conc_317_9;
  wire [7:0] layer4_out_conc_317_8_1;
  wire layer4_out_conc_317_0;
  wire layer4_out_conc_319_9;
  wire [7:0] layer4_out_conc_319_8_1;
  wire layer4_out_conc_319_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_0;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_9;
  wire [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_8_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_0;
  wire [10:0] Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1;
  wire [10:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1;
  wire [10:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire [15:0] Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;
  wire [15:0] Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1;

  wire[15:0] Accum2_1_acc_386_nl;
  wire[21:0] nl_Accum2_1_acc_386_nl;
  wire[14:0] Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_90_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_90_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_91_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_91_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_92_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_92_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_93_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_93_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_94_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_94_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_95_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_95_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_96_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_96_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_97_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_97_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_78_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_78_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_79_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_79_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_74_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_74_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_75_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_75_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_76_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_76_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_77_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_77_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_81_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_81_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_86_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_86_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_87_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_87_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_82_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_82_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_83_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_83_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_84_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_84_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_85_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_85_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_88_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_88_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_89_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_89_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_65_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_65_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_70_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_70_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_71_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_71_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_72_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_72_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_73_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_73_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_66_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_66_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_67_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_67_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_68_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_68_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_69_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_69_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_102_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_102_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_103_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_103_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_104_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_104_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_105_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_105_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_98_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_98_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_99_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_99_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_100_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_100_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_101_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_101_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[15:0] Accum2_1_acc_385_nl;
  wire[20:0] nl_Accum2_1_acc_385_nl;
  wire[14:0] Product1_1_126_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_126_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_123_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_123_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_118_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_118_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_115_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_115_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_122_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_122_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_119_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_119_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_114_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_114_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_111_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_111_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_112_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_112_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_109_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_109_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_389_nl;
  wire[6:0] nl_Accum2_1_acc_389_nl;
  wire[14:0] Product1_1_110_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_110_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_108_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_108_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_127_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_127_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_106_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_106_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_107_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_107_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_128_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_128_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_125_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_125_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_124_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_124_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_121_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_121_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_120_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_120_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_117_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_117_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_116_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_116_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_113_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_113_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[15:0] Accum2_1_acc_259_nl;
  wire[21:0] nl_Accum2_1_acc_259_nl;
  wire[14:0] Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_90_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_90_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_91_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_91_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_92_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_92_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_93_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_93_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_94_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_94_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_95_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_95_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_96_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_96_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_97_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_97_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_78_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_78_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_79_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_79_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_74_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_74_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_75_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_75_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_76_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_76_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_77_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_77_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_80_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_80_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_81_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_81_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_86_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_86_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_87_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_87_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_82_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_82_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_83_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_83_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_84_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_84_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_85_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_85_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_88_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_88_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_89_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_89_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_65_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_65_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_70_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_70_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_71_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_71_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_72_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_72_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_73_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_73_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_66_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_66_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_67_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_67_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_68_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_68_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_69_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_69_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_102_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_102_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_103_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_103_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_104_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_104_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_105_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_105_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_98_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_98_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_99_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_99_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_100_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_100_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_101_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_101_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[15:0] Accum2_1_acc_258_nl;
  wire[20:0] nl_Accum2_1_acc_258_nl;
  wire[14:0] Product1_1_126_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_126_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_123_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_123_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_118_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_118_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_115_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_115_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_122_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_122_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_119_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_119_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_114_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_114_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_111_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_111_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_112_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_112_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_109_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_109_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_388_nl;
  wire[6:0] nl_Accum2_1_acc_388_nl;
  wire[14:0] Product1_1_110_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_110_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_108_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_108_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_127_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_127_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_106_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_106_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_107_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_107_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_128_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_128_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_125_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_125_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_124_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_124_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_121_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_121_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_120_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_120_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_117_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_117_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_116_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_116_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_113_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_113_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[15:0] Accum2_1_acc_132_nl;
  wire[21:0] nl_Accum2_1_acc_132_nl;
  wire[14:0] Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_89_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_89_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_90_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_90_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_91_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_91_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_92_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_92_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_93_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_93_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_94_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_94_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_95_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_95_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_96_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_96_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_77_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_77_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_78_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_78_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_73_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_73_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_74_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_74_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_75_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_75_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_76_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_76_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_79_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_79_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_80_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_80_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_85_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_85_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_86_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_86_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_81_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_81_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_82_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_82_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_83_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_83_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_84_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_84_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_87_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_87_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_88_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_88_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_69_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_69_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_70_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_70_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_71_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_71_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_72_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_72_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_65_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_65_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_66_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_66_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_67_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_67_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_68_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_68_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_101_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_101_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_102_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_102_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_103_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_103_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_104_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_104_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_97_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_97_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_98_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_98_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_99_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_99_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_100_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_100_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[15:0] Accum2_1_acc_131_nl;
  wire[20:0] nl_Accum2_1_acc_131_nl;
  wire[14:0] Product1_1_124_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_124_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_125_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_125_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_116_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_116_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_117_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_117_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_120_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_120_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_121_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_121_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_112_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_112_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_113_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_113_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_110_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_110_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_111_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_111_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_390_nl;
  wire[6:0] nl_Accum2_1_acc_390_nl;
  wire[14:0] Product1_1_108_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_108_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_109_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_109_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_126_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_126_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_105_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_105_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_106_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_106_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_127_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_127_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_128_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_128_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_122_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_122_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_123_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_123_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_118_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_118_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_119_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_119_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_114_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_114_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_115_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_115_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_140_nl;
  wire[17:0] nl_Accum2_acc_140_nl;
  wire[15:0] Accum2_acc_134_nl;
  wire[16:0] nl_Accum2_acc_134_nl;
  wire[19:0] Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_133_nl;
  wire[16:0] nl_Accum2_acc_133_nl;
  wire[19:0] Product1_4_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_132_nl;
  wire[16:0] nl_Accum2_acc_132_nl;
  wire[19:0] Product1_6_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_131_nl;
  wire[16:0] nl_Accum2_acc_131_nl;
  wire[19:0] Product1_8_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_nl;
  wire[16:0] nl_Accum2_acc_nl;
  wire[15:0] Accum2_acc_136_nl;
  wire[16:0] nl_Accum2_acc_136_nl;
  wire[15:0] Accum2_acc_130_nl;
  wire[16:0] nl_Accum2_acc_130_nl;
  wire[19:0] Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_129_nl;
  wire[16:0] nl_Accum2_acc_129_nl;
  wire[19:0] Product1_12_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_139_nl;
  wire[16:0] nl_Accum2_acc_139_nl;
  wire[9:0] Accum2_acc_1792_nl;
  wire[10:0] nl_Accum2_acc_1792_nl;
  wire[19:0] Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_153_nl;
  wire[17:0] nl_Accum2_acc_153_nl;
  wire[15:0] Accum2_acc_147_nl;
  wire[16:0] nl_Accum2_acc_147_nl;
  wire[19:0] Product1_2_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_146_nl;
  wire[16:0] nl_Accum2_acc_146_nl;
  wire[19:0] Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_145_nl;
  wire[16:0] nl_Accum2_acc_145_nl;
  wire[19:0] Product1_6_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_144_nl;
  wire[16:0] nl_Accum2_acc_144_nl;
  wire[19:0] Product1_8_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_152_nl;
  wire[16:0] nl_Accum2_acc_152_nl;
  wire[15:0] Accum2_acc_149_nl;
  wire[16:0] nl_Accum2_acc_149_nl;
  wire[15:0] Accum2_acc_143_nl;
  wire[16:0] nl_Accum2_acc_143_nl;
  wire[19:0] Product1_10_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_142_nl;
  wire[16:0] nl_Accum2_acc_142_nl;
  wire[19:0] Product1_12_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_148_nl;
  wire[16:0] nl_Accum2_acc_148_nl;
  wire[9:0] Accum2_acc_1793_nl;
  wire[10:0] nl_Accum2_acc_1793_nl;
  wire[19:0] Product1_1_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_166_nl;
  wire[17:0] nl_Accum2_acc_166_nl;
  wire[15:0] Accum2_acc_160_nl;
  wire[16:0] nl_Accum2_acc_160_nl;
  wire[19:0] Product1_2_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_159_nl;
  wire[16:0] nl_Accum2_acc_159_nl;
  wire[19:0] Product1_4_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_158_nl;
  wire[16:0] nl_Accum2_acc_158_nl;
  wire[19:0] Product1_6_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_157_nl;
  wire[16:0] nl_Accum2_acc_157_nl;
  wire[19:0] Product1_8_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_165_nl;
  wire[16:0] nl_Accum2_acc_165_nl;
  wire[15:0] Accum2_acc_162_nl;
  wire[16:0] nl_Accum2_acc_162_nl;
  wire[15:0] Accum2_acc_156_nl;
  wire[16:0] nl_Accum2_acc_156_nl;
  wire[19:0] Product1_10_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_155_nl;
  wire[16:0] nl_Accum2_acc_155_nl;
  wire[19:0] Product1_12_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_161_nl;
  wire[16:0] nl_Accum2_acc_161_nl;
  wire[9:0] Accum2_acc_1794_nl;
  wire[10:0] nl_Accum2_acc_1794_nl;
  wire[19:0] Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_179_nl;
  wire[17:0] nl_Accum2_acc_179_nl;
  wire[15:0] Accum2_acc_173_nl;
  wire[16:0] nl_Accum2_acc_173_nl;
  wire[19:0] Product1_2_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_172_nl;
  wire[16:0] nl_Accum2_acc_172_nl;
  wire[19:0] Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_171_nl;
  wire[16:0] nl_Accum2_acc_171_nl;
  wire[19:0] Product1_6_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_170_nl;
  wire[16:0] nl_Accum2_acc_170_nl;
  wire[19:0] Product1_8_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_178_nl;
  wire[16:0] nl_Accum2_acc_178_nl;
  wire[15:0] Accum2_acc_175_nl;
  wire[16:0] nl_Accum2_acc_175_nl;
  wire[15:0] Accum2_acc_169_nl;
  wire[16:0] nl_Accum2_acc_169_nl;
  wire[19:0] Product1_10_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_168_nl;
  wire[16:0] nl_Accum2_acc_168_nl;
  wire[19:0] Product1_12_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_174_nl;
  wire[16:0] nl_Accum2_acc_174_nl;
  wire[9:0] Accum2_acc_1795_nl;
  wire[10:0] nl_Accum2_acc_1795_nl;
  wire[19:0] Product1_1_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_192_nl;
  wire[17:0] nl_Accum2_acc_192_nl;
  wire[15:0] Accum2_acc_186_nl;
  wire[16:0] nl_Accum2_acc_186_nl;
  wire[19:0] Product1_2_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_185_nl;
  wire[16:0] nl_Accum2_acc_185_nl;
  wire[19:0] Product1_4_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_184_nl;
  wire[16:0] nl_Accum2_acc_184_nl;
  wire[19:0] Product1_6_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_183_nl;
  wire[16:0] nl_Accum2_acc_183_nl;
  wire[19:0] Product1_8_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_191_nl;
  wire[16:0] nl_Accum2_acc_191_nl;
  wire[15:0] Accum2_acc_188_nl;
  wire[16:0] nl_Accum2_acc_188_nl;
  wire[15:0] Accum2_acc_182_nl;
  wire[16:0] nl_Accum2_acc_182_nl;
  wire[19:0] Product1_10_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_181_nl;
  wire[16:0] nl_Accum2_acc_181_nl;
  wire[19:0] Product1_12_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_187_nl;
  wire[16:0] nl_Accum2_acc_187_nl;
  wire[9:0] Accum2_acc_1796_nl;
  wire[10:0] nl_Accum2_acc_1796_nl;
  wire[19:0] Product1_1_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_205_nl;
  wire[17:0] nl_Accum2_acc_205_nl;
  wire[15:0] Accum2_acc_199_nl;
  wire[16:0] nl_Accum2_acc_199_nl;
  wire[19:0] Product1_2_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_198_nl;
  wire[16:0] nl_Accum2_acc_198_nl;
  wire[19:0] Product1_4_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_197_nl;
  wire[16:0] nl_Accum2_acc_197_nl;
  wire[19:0] Product1_6_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_196_nl;
  wire[16:0] nl_Accum2_acc_196_nl;
  wire[19:0] Product1_8_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_204_nl;
  wire[16:0] nl_Accum2_acc_204_nl;
  wire[15:0] Accum2_acc_201_nl;
  wire[16:0] nl_Accum2_acc_201_nl;
  wire[15:0] Accum2_acc_195_nl;
  wire[16:0] nl_Accum2_acc_195_nl;
  wire[19:0] Product1_10_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_194_nl;
  wire[16:0] nl_Accum2_acc_194_nl;
  wire[19:0] Product1_12_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_200_nl;
  wire[16:0] nl_Accum2_acc_200_nl;
  wire[9:0] Accum2_acc_1797_nl;
  wire[10:0] nl_Accum2_acc_1797_nl;
  wire[19:0] Product1_1_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_218_nl;
  wire[17:0] nl_Accum2_acc_218_nl;
  wire[15:0] Accum2_acc_212_nl;
  wire[16:0] nl_Accum2_acc_212_nl;
  wire[19:0] Product1_2_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_211_nl;
  wire[16:0] nl_Accum2_acc_211_nl;
  wire[19:0] Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_210_nl;
  wire[16:0] nl_Accum2_acc_210_nl;
  wire[19:0] Product1_6_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_209_nl;
  wire[16:0] nl_Accum2_acc_209_nl;
  wire[19:0] Product1_8_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_217_nl;
  wire[16:0] nl_Accum2_acc_217_nl;
  wire[15:0] Accum2_acc_214_nl;
  wire[16:0] nl_Accum2_acc_214_nl;
  wire[15:0] Accum2_acc_208_nl;
  wire[16:0] nl_Accum2_acc_208_nl;
  wire[19:0] Product1_10_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_207_nl;
  wire[16:0] nl_Accum2_acc_207_nl;
  wire[19:0] Product1_12_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_213_nl;
  wire[16:0] nl_Accum2_acc_213_nl;
  wire[9:0] Accum2_acc_1798_nl;
  wire[10:0] nl_Accum2_acc_1798_nl;
  wire[19:0] Product1_1_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_231_nl;
  wire[17:0] nl_Accum2_acc_231_nl;
  wire[15:0] Accum2_acc_225_nl;
  wire[16:0] nl_Accum2_acc_225_nl;
  wire[19:0] Product1_2_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_224_nl;
  wire[16:0] nl_Accum2_acc_224_nl;
  wire[19:0] Product1_4_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_223_nl;
  wire[16:0] nl_Accum2_acc_223_nl;
  wire[19:0] Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_222_nl;
  wire[16:0] nl_Accum2_acc_222_nl;
  wire[19:0] Product1_8_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_230_nl;
  wire[16:0] nl_Accum2_acc_230_nl;
  wire[15:0] Accum2_acc_227_nl;
  wire[16:0] nl_Accum2_acc_227_nl;
  wire[15:0] Accum2_acc_221_nl;
  wire[16:0] nl_Accum2_acc_221_nl;
  wire[19:0] Product1_10_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_220_nl;
  wire[16:0] nl_Accum2_acc_220_nl;
  wire[19:0] Product1_12_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_226_nl;
  wire[16:0] nl_Accum2_acc_226_nl;
  wire[9:0] Accum2_acc_1799_nl;
  wire[10:0] nl_Accum2_acc_1799_nl;
  wire[19:0] Product1_1_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_244_nl;
  wire[17:0] nl_Accum2_acc_244_nl;
  wire[15:0] Accum2_acc_238_nl;
  wire[16:0] nl_Accum2_acc_238_nl;
  wire[19:0] Product1_2_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_237_nl;
  wire[16:0] nl_Accum2_acc_237_nl;
  wire[19:0] Product1_4_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_236_nl;
  wire[16:0] nl_Accum2_acc_236_nl;
  wire[19:0] Product1_6_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_235_nl;
  wire[16:0] nl_Accum2_acc_235_nl;
  wire[19:0] Product1_8_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_243_nl;
  wire[16:0] nl_Accum2_acc_243_nl;
  wire[15:0] Accum2_acc_240_nl;
  wire[16:0] nl_Accum2_acc_240_nl;
  wire[15:0] Accum2_acc_234_nl;
  wire[16:0] nl_Accum2_acc_234_nl;
  wire[19:0] Product1_10_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_233_nl;
  wire[16:0] nl_Accum2_acc_233_nl;
  wire[19:0] Product1_12_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_239_nl;
  wire[16:0] nl_Accum2_acc_239_nl;
  wire[9:0] Accum2_acc_1800_nl;
  wire[10:0] nl_Accum2_acc_1800_nl;
  wire[19:0] Product1_1_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_257_nl;
  wire[17:0] nl_Accum2_acc_257_nl;
  wire[15:0] Accum2_acc_251_nl;
  wire[16:0] nl_Accum2_acc_251_nl;
  wire[19:0] Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_250_nl;
  wire[16:0] nl_Accum2_acc_250_nl;
  wire[19:0] Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_249_nl;
  wire[16:0] nl_Accum2_acc_249_nl;
  wire[19:0] Product1_6_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_248_nl;
  wire[16:0] nl_Accum2_acc_248_nl;
  wire[19:0] Product1_8_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_256_nl;
  wire[16:0] nl_Accum2_acc_256_nl;
  wire[15:0] Accum2_acc_253_nl;
  wire[16:0] nl_Accum2_acc_253_nl;
  wire[15:0] Accum2_acc_247_nl;
  wire[16:0] nl_Accum2_acc_247_nl;
  wire[19:0] Product1_10_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_246_nl;
  wire[16:0] nl_Accum2_acc_246_nl;
  wire[19:0] Product1_12_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_252_nl;
  wire[16:0] nl_Accum2_acc_252_nl;
  wire[9:0] Accum2_acc_1801_nl;
  wire[10:0] nl_Accum2_acc_1801_nl;
  wire[19:0] Product1_1_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_270_nl;
  wire[17:0] nl_Accum2_acc_270_nl;
  wire[15:0] Accum2_acc_264_nl;
  wire[16:0] nl_Accum2_acc_264_nl;
  wire[19:0] Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_263_nl;
  wire[16:0] nl_Accum2_acc_263_nl;
  wire[19:0] Product1_4_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_262_nl;
  wire[16:0] nl_Accum2_acc_262_nl;
  wire[19:0] Product1_6_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_261_nl;
  wire[16:0] nl_Accum2_acc_261_nl;
  wire[19:0] Product1_8_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_269_nl;
  wire[16:0] nl_Accum2_acc_269_nl;
  wire[15:0] Accum2_acc_266_nl;
  wire[16:0] nl_Accum2_acc_266_nl;
  wire[15:0] Accum2_acc_260_nl;
  wire[16:0] nl_Accum2_acc_260_nl;
  wire[19:0] Product1_10_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_259_nl;
  wire[16:0] nl_Accum2_acc_259_nl;
  wire[19:0] Product1_12_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_265_nl;
  wire[16:0] nl_Accum2_acc_265_nl;
  wire[9:0] Accum2_acc_1802_nl;
  wire[10:0] nl_Accum2_acc_1802_nl;
  wire[19:0] Product1_1_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_283_nl;
  wire[17:0] nl_Accum2_acc_283_nl;
  wire[15:0] Accum2_acc_277_nl;
  wire[16:0] nl_Accum2_acc_277_nl;
  wire[19:0] Product1_2_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_276_nl;
  wire[16:0] nl_Accum2_acc_276_nl;
  wire[19:0] Product1_4_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_275_nl;
  wire[16:0] nl_Accum2_acc_275_nl;
  wire[19:0] Product1_6_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_274_nl;
  wire[16:0] nl_Accum2_acc_274_nl;
  wire[19:0] Product1_8_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_282_nl;
  wire[16:0] nl_Accum2_acc_282_nl;
  wire[15:0] Accum2_acc_279_nl;
  wire[16:0] nl_Accum2_acc_279_nl;
  wire[15:0] Accum2_acc_273_nl;
  wire[16:0] nl_Accum2_acc_273_nl;
  wire[19:0] Product1_10_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_272_nl;
  wire[16:0] nl_Accum2_acc_272_nl;
  wire[19:0] Product1_12_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_278_nl;
  wire[16:0] nl_Accum2_acc_278_nl;
  wire[9:0] Accum2_acc_1803_nl;
  wire[10:0] nl_Accum2_acc_1803_nl;
  wire[19:0] Product1_1_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_296_nl;
  wire[17:0] nl_Accum2_acc_296_nl;
  wire[15:0] Accum2_acc_290_nl;
  wire[16:0] nl_Accum2_acc_290_nl;
  wire[19:0] Product1_2_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_289_nl;
  wire[16:0] nl_Accum2_acc_289_nl;
  wire[19:0] Product1_4_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_288_nl;
  wire[16:0] nl_Accum2_acc_288_nl;
  wire[19:0] Product1_6_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_287_nl;
  wire[16:0] nl_Accum2_acc_287_nl;
  wire[19:0] Product1_8_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_295_nl;
  wire[16:0] nl_Accum2_acc_295_nl;
  wire[15:0] Accum2_acc_292_nl;
  wire[16:0] nl_Accum2_acc_292_nl;
  wire[15:0] Accum2_acc_286_nl;
  wire[16:0] nl_Accum2_acc_286_nl;
  wire[19:0] Product1_10_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_285_nl;
  wire[16:0] nl_Accum2_acc_285_nl;
  wire[19:0] Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_291_nl;
  wire[16:0] nl_Accum2_acc_291_nl;
  wire[9:0] Accum2_acc_1804_nl;
  wire[10:0] nl_Accum2_acc_1804_nl;
  wire[19:0] Product1_1_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_309_nl;
  wire[17:0] nl_Accum2_acc_309_nl;
  wire[15:0] Accum2_acc_303_nl;
  wire[16:0] nl_Accum2_acc_303_nl;
  wire[19:0] Product1_2_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_302_nl;
  wire[16:0] nl_Accum2_acc_302_nl;
  wire[19:0] Product1_4_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_301_nl;
  wire[16:0] nl_Accum2_acc_301_nl;
  wire[19:0] Product1_6_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_300_nl;
  wire[16:0] nl_Accum2_acc_300_nl;
  wire[19:0] Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_308_nl;
  wire[16:0] nl_Accum2_acc_308_nl;
  wire[15:0] Accum2_acc_305_nl;
  wire[16:0] nl_Accum2_acc_305_nl;
  wire[15:0] Accum2_acc_299_nl;
  wire[16:0] nl_Accum2_acc_299_nl;
  wire[19:0] Product1_10_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_298_nl;
  wire[16:0] nl_Accum2_acc_298_nl;
  wire[19:0] Product1_12_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_304_nl;
  wire[16:0] nl_Accum2_acc_304_nl;
  wire[9:0] Accum2_acc_1805_nl;
  wire[10:0] nl_Accum2_acc_1805_nl;
  wire[19:0] Product1_1_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_322_nl;
  wire[17:0] nl_Accum2_acc_322_nl;
  wire[15:0] Accum2_acc_316_nl;
  wire[16:0] nl_Accum2_acc_316_nl;
  wire[19:0] Product1_2_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_315_nl;
  wire[16:0] nl_Accum2_acc_315_nl;
  wire[19:0] Product1_4_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_314_nl;
  wire[16:0] nl_Accum2_acc_314_nl;
  wire[19:0] Product1_6_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_313_nl;
  wire[16:0] nl_Accum2_acc_313_nl;
  wire[19:0] Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_321_nl;
  wire[16:0] nl_Accum2_acc_321_nl;
  wire[15:0] Accum2_acc_318_nl;
  wire[16:0] nl_Accum2_acc_318_nl;
  wire[15:0] Accum2_acc_312_nl;
  wire[16:0] nl_Accum2_acc_312_nl;
  wire[19:0] Product1_10_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_311_nl;
  wire[16:0] nl_Accum2_acc_311_nl;
  wire[19:0] Product1_12_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_317_nl;
  wire[16:0] nl_Accum2_acc_317_nl;
  wire[9:0] Accum2_acc_1806_nl;
  wire[10:0] nl_Accum2_acc_1806_nl;
  wire[19:0] Product1_1_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_335_nl;
  wire[17:0] nl_Accum2_acc_335_nl;
  wire[15:0] Accum2_acc_329_nl;
  wire[16:0] nl_Accum2_acc_329_nl;
  wire[19:0] Product1_2_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_328_nl;
  wire[16:0] nl_Accum2_acc_328_nl;
  wire[19:0] Product1_4_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_327_nl;
  wire[16:0] nl_Accum2_acc_327_nl;
  wire[19:0] Product1_6_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_326_nl;
  wire[16:0] nl_Accum2_acc_326_nl;
  wire[19:0] Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_334_nl;
  wire[16:0] nl_Accum2_acc_334_nl;
  wire[15:0] Accum2_acc_331_nl;
  wire[16:0] nl_Accum2_acc_331_nl;
  wire[15:0] Accum2_acc_325_nl;
  wire[16:0] nl_Accum2_acc_325_nl;
  wire[19:0] Product1_10_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_324_nl;
  wire[16:0] nl_Accum2_acc_324_nl;
  wire[19:0] Product1_12_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_330_nl;
  wire[16:0] nl_Accum2_acc_330_nl;
  wire[9:0] Accum2_acc_1807_nl;
  wire[10:0] nl_Accum2_acc_1807_nl;
  wire[19:0] Product1_1_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_348_nl;
  wire[17:0] nl_Accum2_acc_348_nl;
  wire[15:0] Accum2_acc_342_nl;
  wire[16:0] nl_Accum2_acc_342_nl;
  wire[19:0] Product1_2_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_341_nl;
  wire[16:0] nl_Accum2_acc_341_nl;
  wire[19:0] Product1_4_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_340_nl;
  wire[16:0] nl_Accum2_acc_340_nl;
  wire[19:0] Product1_6_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_339_nl;
  wire[16:0] nl_Accum2_acc_339_nl;
  wire[19:0] Product1_8_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_347_nl;
  wire[16:0] nl_Accum2_acc_347_nl;
  wire[15:0] Accum2_acc_344_nl;
  wire[16:0] nl_Accum2_acc_344_nl;
  wire[15:0] Accum2_acc_338_nl;
  wire[16:0] nl_Accum2_acc_338_nl;
  wire[19:0] Product1_10_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_337_nl;
  wire[16:0] nl_Accum2_acc_337_nl;
  wire[19:0] Product1_12_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_343_nl;
  wire[16:0] nl_Accum2_acc_343_nl;
  wire[9:0] Accum2_acc_1808_nl;
  wire[10:0] nl_Accum2_acc_1808_nl;
  wire[19:0] Product1_1_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_361_nl;
  wire[17:0] nl_Accum2_acc_361_nl;
  wire[15:0] Accum2_acc_355_nl;
  wire[16:0] nl_Accum2_acc_355_nl;
  wire[19:0] Product1_2_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_354_nl;
  wire[16:0] nl_Accum2_acc_354_nl;
  wire[19:0] Product1_4_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_353_nl;
  wire[16:0] nl_Accum2_acc_353_nl;
  wire[19:0] Product1_6_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_352_nl;
  wire[16:0] nl_Accum2_acc_352_nl;
  wire[19:0] Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_360_nl;
  wire[16:0] nl_Accum2_acc_360_nl;
  wire[15:0] Accum2_acc_357_nl;
  wire[16:0] nl_Accum2_acc_357_nl;
  wire[15:0] Accum2_acc_351_nl;
  wire[16:0] nl_Accum2_acc_351_nl;
  wire[19:0] Product1_10_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_350_nl;
  wire[16:0] nl_Accum2_acc_350_nl;
  wire[19:0] Product1_12_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_356_nl;
  wire[16:0] nl_Accum2_acc_356_nl;
  wire[9:0] Accum2_acc_1809_nl;
  wire[10:0] nl_Accum2_acc_1809_nl;
  wire[19:0] Product1_1_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_374_nl;
  wire[17:0] nl_Accum2_acc_374_nl;
  wire[15:0] Accum2_acc_368_nl;
  wire[16:0] nl_Accum2_acc_368_nl;
  wire[19:0] Product1_2_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_367_nl;
  wire[16:0] nl_Accum2_acc_367_nl;
  wire[19:0] Product1_4_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_366_nl;
  wire[16:0] nl_Accum2_acc_366_nl;
  wire[19:0] Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_365_nl;
  wire[16:0] nl_Accum2_acc_365_nl;
  wire[19:0] Product1_8_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_373_nl;
  wire[16:0] nl_Accum2_acc_373_nl;
  wire[15:0] Accum2_acc_370_nl;
  wire[16:0] nl_Accum2_acc_370_nl;
  wire[15:0] Accum2_acc_364_nl;
  wire[16:0] nl_Accum2_acc_364_nl;
  wire[19:0] Product1_10_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_363_nl;
  wire[16:0] nl_Accum2_acc_363_nl;
  wire[19:0] Product1_12_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_369_nl;
  wire[16:0] nl_Accum2_acc_369_nl;
  wire[9:0] Accum2_acc_1810_nl;
  wire[10:0] nl_Accum2_acc_1810_nl;
  wire[19:0] Product1_1_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_387_nl;
  wire[17:0] nl_Accum2_acc_387_nl;
  wire[15:0] Accum2_acc_381_nl;
  wire[16:0] nl_Accum2_acc_381_nl;
  wire[19:0] Product1_2_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_380_nl;
  wire[16:0] nl_Accum2_acc_380_nl;
  wire[19:0] Product1_4_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_379_nl;
  wire[16:0] nl_Accum2_acc_379_nl;
  wire[19:0] Product1_6_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_378_nl;
  wire[16:0] nl_Accum2_acc_378_nl;
  wire[19:0] Product1_8_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_386_nl;
  wire[16:0] nl_Accum2_acc_386_nl;
  wire[15:0] Accum2_acc_383_nl;
  wire[16:0] nl_Accum2_acc_383_nl;
  wire[15:0] Accum2_acc_377_nl;
  wire[16:0] nl_Accum2_acc_377_nl;
  wire[19:0] Product1_10_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_376_nl;
  wire[16:0] nl_Accum2_acc_376_nl;
  wire[19:0] Product1_12_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_382_nl;
  wire[16:0] nl_Accum2_acc_382_nl;
  wire[9:0] Accum2_acc_1811_nl;
  wire[10:0] nl_Accum2_acc_1811_nl;
  wire[19:0] Product1_1_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_400_nl;
  wire[17:0] nl_Accum2_acc_400_nl;
  wire[15:0] Accum2_acc_394_nl;
  wire[16:0] nl_Accum2_acc_394_nl;
  wire[19:0] Product1_2_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_393_nl;
  wire[16:0] nl_Accum2_acc_393_nl;
  wire[19:0] Product1_4_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_392_nl;
  wire[16:0] nl_Accum2_acc_392_nl;
  wire[19:0] Product1_6_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_391_nl;
  wire[16:0] nl_Accum2_acc_391_nl;
  wire[19:0] Product1_8_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_399_nl;
  wire[16:0] nl_Accum2_acc_399_nl;
  wire[15:0] Accum2_acc_396_nl;
  wire[16:0] nl_Accum2_acc_396_nl;
  wire[15:0] Accum2_acc_390_nl;
  wire[16:0] nl_Accum2_acc_390_nl;
  wire[19:0] Product1_10_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_389_nl;
  wire[16:0] nl_Accum2_acc_389_nl;
  wire[19:0] Product1_12_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_395_nl;
  wire[16:0] nl_Accum2_acc_395_nl;
  wire[9:0] Accum2_acc_1812_nl;
  wire[10:0] nl_Accum2_acc_1812_nl;
  wire[19:0] Product1_1_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_413_nl;
  wire[17:0] nl_Accum2_acc_413_nl;
  wire[15:0] Accum2_acc_407_nl;
  wire[16:0] nl_Accum2_acc_407_nl;
  wire[19:0] Product1_2_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_406_nl;
  wire[16:0] nl_Accum2_acc_406_nl;
  wire[19:0] Product1_4_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_405_nl;
  wire[16:0] nl_Accum2_acc_405_nl;
  wire[19:0] Product1_6_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_404_nl;
  wire[16:0] nl_Accum2_acc_404_nl;
  wire[19:0] Product1_8_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_412_nl;
  wire[16:0] nl_Accum2_acc_412_nl;
  wire[15:0] Accum2_acc_409_nl;
  wire[16:0] nl_Accum2_acc_409_nl;
  wire[15:0] Accum2_acc_403_nl;
  wire[16:0] nl_Accum2_acc_403_nl;
  wire[19:0] Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_402_nl;
  wire[16:0] nl_Accum2_acc_402_nl;
  wire[19:0] Product1_12_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_408_nl;
  wire[16:0] nl_Accum2_acc_408_nl;
  wire[9:0] Accum2_acc_1813_nl;
  wire[10:0] nl_Accum2_acc_1813_nl;
  wire[19:0] Product1_1_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_426_nl;
  wire[17:0] nl_Accum2_acc_426_nl;
  wire[15:0] Accum2_acc_420_nl;
  wire[16:0] nl_Accum2_acc_420_nl;
  wire[19:0] Product1_2_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_419_nl;
  wire[16:0] nl_Accum2_acc_419_nl;
  wire[19:0] Product1_4_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_418_nl;
  wire[16:0] nl_Accum2_acc_418_nl;
  wire[19:0] Product1_6_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_417_nl;
  wire[16:0] nl_Accum2_acc_417_nl;
  wire[19:0] Product1_8_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_425_nl;
  wire[16:0] nl_Accum2_acc_425_nl;
  wire[15:0] Accum2_acc_422_nl;
  wire[16:0] nl_Accum2_acc_422_nl;
  wire[15:0] Accum2_acc_416_nl;
  wire[16:0] nl_Accum2_acc_416_nl;
  wire[19:0] Product1_10_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_415_nl;
  wire[16:0] nl_Accum2_acc_415_nl;
  wire[19:0] Product1_12_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_421_nl;
  wire[16:0] nl_Accum2_acc_421_nl;
  wire[9:0] Accum2_acc_1814_nl;
  wire[10:0] nl_Accum2_acc_1814_nl;
  wire[19:0] Product1_1_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_439_nl;
  wire[17:0] nl_Accum2_acc_439_nl;
  wire[15:0] Accum2_acc_433_nl;
  wire[16:0] nl_Accum2_acc_433_nl;
  wire[19:0] Product1_2_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_432_nl;
  wire[16:0] nl_Accum2_acc_432_nl;
  wire[19:0] Product1_4_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_431_nl;
  wire[16:0] nl_Accum2_acc_431_nl;
  wire[19:0] Product1_6_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_430_nl;
  wire[16:0] nl_Accum2_acc_430_nl;
  wire[19:0] Product1_8_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_438_nl;
  wire[16:0] nl_Accum2_acc_438_nl;
  wire[15:0] Accum2_acc_435_nl;
  wire[16:0] nl_Accum2_acc_435_nl;
  wire[15:0] Accum2_acc_429_nl;
  wire[16:0] nl_Accum2_acc_429_nl;
  wire[19:0] Product1_10_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_428_nl;
  wire[16:0] nl_Accum2_acc_428_nl;
  wire[19:0] Product1_12_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_434_nl;
  wire[16:0] nl_Accum2_acc_434_nl;
  wire[9:0] Accum2_acc_1815_nl;
  wire[10:0] nl_Accum2_acc_1815_nl;
  wire[19:0] Product1_1_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_452_nl;
  wire[17:0] nl_Accum2_acc_452_nl;
  wire[15:0] Accum2_acc_446_nl;
  wire[16:0] nl_Accum2_acc_446_nl;
  wire[19:0] Product1_2_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_445_nl;
  wire[16:0] nl_Accum2_acc_445_nl;
  wire[19:0] Product1_4_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_444_nl;
  wire[16:0] nl_Accum2_acc_444_nl;
  wire[19:0] Product1_6_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_443_nl;
  wire[16:0] nl_Accum2_acc_443_nl;
  wire[19:0] Product1_8_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_451_nl;
  wire[16:0] nl_Accum2_acc_451_nl;
  wire[15:0] Accum2_acc_448_nl;
  wire[16:0] nl_Accum2_acc_448_nl;
  wire[15:0] Accum2_acc_442_nl;
  wire[16:0] nl_Accum2_acc_442_nl;
  wire[19:0] Product1_10_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_441_nl;
  wire[16:0] nl_Accum2_acc_441_nl;
  wire[19:0] Product1_12_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_447_nl;
  wire[16:0] nl_Accum2_acc_447_nl;
  wire[9:0] Accum2_acc_1816_nl;
  wire[10:0] nl_Accum2_acc_1816_nl;
  wire[19:0] Product1_1_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_465_nl;
  wire[17:0] nl_Accum2_acc_465_nl;
  wire[15:0] Accum2_acc_459_nl;
  wire[16:0] nl_Accum2_acc_459_nl;
  wire[19:0] Product1_2_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_458_nl;
  wire[16:0] nl_Accum2_acc_458_nl;
  wire[19:0] Product1_4_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_457_nl;
  wire[16:0] nl_Accum2_acc_457_nl;
  wire[19:0] Product1_6_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_456_nl;
  wire[16:0] nl_Accum2_acc_456_nl;
  wire[19:0] Product1_8_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_464_nl;
  wire[16:0] nl_Accum2_acc_464_nl;
  wire[15:0] Accum2_acc_461_nl;
  wire[16:0] nl_Accum2_acc_461_nl;
  wire[15:0] Accum2_acc_455_nl;
  wire[16:0] nl_Accum2_acc_455_nl;
  wire[19:0] Product1_10_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_454_nl;
  wire[16:0] nl_Accum2_acc_454_nl;
  wire[19:0] Product1_12_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_460_nl;
  wire[16:0] nl_Accum2_acc_460_nl;
  wire[9:0] Accum2_acc_1817_nl;
  wire[10:0] nl_Accum2_acc_1817_nl;
  wire[19:0] Product1_1_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_478_nl;
  wire[17:0] nl_Accum2_acc_478_nl;
  wire[15:0] Accum2_acc_472_nl;
  wire[16:0] nl_Accum2_acc_472_nl;
  wire[19:0] Product1_2_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_471_nl;
  wire[16:0] nl_Accum2_acc_471_nl;
  wire[19:0] Product1_4_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_470_nl;
  wire[16:0] nl_Accum2_acc_470_nl;
  wire[19:0] Product1_6_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_469_nl;
  wire[16:0] nl_Accum2_acc_469_nl;
  wire[19:0] Product1_8_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_477_nl;
  wire[16:0] nl_Accum2_acc_477_nl;
  wire[15:0] Accum2_acc_474_nl;
  wire[16:0] nl_Accum2_acc_474_nl;
  wire[15:0] Accum2_acc_468_nl;
  wire[16:0] nl_Accum2_acc_468_nl;
  wire[19:0] Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_467_nl;
  wire[16:0] nl_Accum2_acc_467_nl;
  wire[19:0] Product1_12_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_473_nl;
  wire[16:0] nl_Accum2_acc_473_nl;
  wire[9:0] Accum2_acc_1818_nl;
  wire[10:0] nl_Accum2_acc_1818_nl;
  wire[19:0] Product1_1_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_491_nl;
  wire[17:0] nl_Accum2_acc_491_nl;
  wire[15:0] Accum2_acc_485_nl;
  wire[16:0] nl_Accum2_acc_485_nl;
  wire[19:0] Product1_2_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_484_nl;
  wire[16:0] nl_Accum2_acc_484_nl;
  wire[19:0] Product1_4_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_483_nl;
  wire[16:0] nl_Accum2_acc_483_nl;
  wire[19:0] Product1_6_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_482_nl;
  wire[16:0] nl_Accum2_acc_482_nl;
  wire[19:0] Product1_8_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_490_nl;
  wire[16:0] nl_Accum2_acc_490_nl;
  wire[15:0] Accum2_acc_487_nl;
  wire[16:0] nl_Accum2_acc_487_nl;
  wire[15:0] Accum2_acc_481_nl;
  wire[16:0] nl_Accum2_acc_481_nl;
  wire[19:0] Product1_10_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_480_nl;
  wire[16:0] nl_Accum2_acc_480_nl;
  wire[19:0] Product1_12_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_486_nl;
  wire[16:0] nl_Accum2_acc_486_nl;
  wire[9:0] Accum2_acc_1819_nl;
  wire[10:0] nl_Accum2_acc_1819_nl;
  wire[19:0] Product1_1_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_504_nl;
  wire[17:0] nl_Accum2_acc_504_nl;
  wire[15:0] Accum2_acc_498_nl;
  wire[16:0] nl_Accum2_acc_498_nl;
  wire[19:0] Product1_2_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_497_nl;
  wire[16:0] nl_Accum2_acc_497_nl;
  wire[19:0] Product1_4_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_496_nl;
  wire[16:0] nl_Accum2_acc_496_nl;
  wire[19:0] Product1_6_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_495_nl;
  wire[16:0] nl_Accum2_acc_495_nl;
  wire[19:0] Product1_8_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_503_nl;
  wire[16:0] nl_Accum2_acc_503_nl;
  wire[15:0] Accum2_acc_500_nl;
  wire[16:0] nl_Accum2_acc_500_nl;
  wire[15:0] Accum2_acc_494_nl;
  wire[16:0] nl_Accum2_acc_494_nl;
  wire[19:0] Product1_10_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_493_nl;
  wire[16:0] nl_Accum2_acc_493_nl;
  wire[19:0] Product1_12_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_499_nl;
  wire[16:0] nl_Accum2_acc_499_nl;
  wire[9:0] Accum2_acc_1820_nl;
  wire[10:0] nl_Accum2_acc_1820_nl;
  wire[19:0] Product1_1_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_517_nl;
  wire[17:0] nl_Accum2_acc_517_nl;
  wire[15:0] Accum2_acc_511_nl;
  wire[16:0] nl_Accum2_acc_511_nl;
  wire[19:0] Product1_2_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_510_nl;
  wire[16:0] nl_Accum2_acc_510_nl;
  wire[19:0] Product1_4_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_509_nl;
  wire[16:0] nl_Accum2_acc_509_nl;
  wire[19:0] Product1_6_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_508_nl;
  wire[16:0] nl_Accum2_acc_508_nl;
  wire[19:0] Product1_8_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_516_nl;
  wire[16:0] nl_Accum2_acc_516_nl;
  wire[15:0] Accum2_acc_513_nl;
  wire[16:0] nl_Accum2_acc_513_nl;
  wire[15:0] Accum2_acc_507_nl;
  wire[16:0] nl_Accum2_acc_507_nl;
  wire[19:0] Product1_10_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_506_nl;
  wire[16:0] nl_Accum2_acc_506_nl;
  wire[19:0] Product1_12_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_512_nl;
  wire[16:0] nl_Accum2_acc_512_nl;
  wire[9:0] Accum2_acc_1821_nl;
  wire[10:0] nl_Accum2_acc_1821_nl;
  wire[19:0] Product1_1_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_530_nl;
  wire[17:0] nl_Accum2_acc_530_nl;
  wire[15:0] Accum2_acc_524_nl;
  wire[16:0] nl_Accum2_acc_524_nl;
  wire[19:0] Product1_2_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_523_nl;
  wire[16:0] nl_Accum2_acc_523_nl;
  wire[19:0] Product1_4_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_522_nl;
  wire[16:0] nl_Accum2_acc_522_nl;
  wire[19:0] Product1_6_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_521_nl;
  wire[16:0] nl_Accum2_acc_521_nl;
  wire[19:0] Product1_8_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_529_nl;
  wire[16:0] nl_Accum2_acc_529_nl;
  wire[15:0] Accum2_acc_526_nl;
  wire[16:0] nl_Accum2_acc_526_nl;
  wire[15:0] Accum2_acc_520_nl;
  wire[16:0] nl_Accum2_acc_520_nl;
  wire[19:0] Product1_10_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_519_nl;
  wire[16:0] nl_Accum2_acc_519_nl;
  wire[19:0] Product1_12_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_525_nl;
  wire[16:0] nl_Accum2_acc_525_nl;
  wire[9:0] Accum2_acc_1822_nl;
  wire[10:0] nl_Accum2_acc_1822_nl;
  wire[19:0] Product1_1_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_543_nl;
  wire[17:0] nl_Accum2_acc_543_nl;
  wire[15:0] Accum2_acc_537_nl;
  wire[16:0] nl_Accum2_acc_537_nl;
  wire[19:0] Product1_2_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_536_nl;
  wire[16:0] nl_Accum2_acc_536_nl;
  wire[19:0] Product1_4_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_535_nl;
  wire[16:0] nl_Accum2_acc_535_nl;
  wire[19:0] Product1_6_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_534_nl;
  wire[16:0] nl_Accum2_acc_534_nl;
  wire[19:0] Product1_8_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_542_nl;
  wire[16:0] nl_Accum2_acc_542_nl;
  wire[15:0] Accum2_acc_539_nl;
  wire[16:0] nl_Accum2_acc_539_nl;
  wire[15:0] Accum2_acc_533_nl;
  wire[16:0] nl_Accum2_acc_533_nl;
  wire[19:0] Product1_10_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_532_nl;
  wire[16:0] nl_Accum2_acc_532_nl;
  wire[19:0] Product1_12_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_538_nl;
  wire[16:0] nl_Accum2_acc_538_nl;
  wire[9:0] Accum2_acc_1823_nl;
  wire[10:0] nl_Accum2_acc_1823_nl;
  wire[19:0] Product1_1_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_556_nl;
  wire[17:0] nl_Accum2_acc_556_nl;
  wire[15:0] Accum2_acc_550_nl;
  wire[16:0] nl_Accum2_acc_550_nl;
  wire[19:0] Product1_2_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_549_nl;
  wire[16:0] nl_Accum2_acc_549_nl;
  wire[19:0] Product1_4_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_548_nl;
  wire[16:0] nl_Accum2_acc_548_nl;
  wire[19:0] Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_547_nl;
  wire[16:0] nl_Accum2_acc_547_nl;
  wire[19:0] Product1_8_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_555_nl;
  wire[16:0] nl_Accum2_acc_555_nl;
  wire[15:0] Accum2_acc_552_nl;
  wire[16:0] nl_Accum2_acc_552_nl;
  wire[15:0] Accum2_acc_546_nl;
  wire[16:0] nl_Accum2_acc_546_nl;
  wire[19:0] Product1_10_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_545_nl;
  wire[16:0] nl_Accum2_acc_545_nl;
  wire[19:0] Product1_12_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_551_nl;
  wire[16:0] nl_Accum2_acc_551_nl;
  wire[9:0] Accum2_acc_1824_nl;
  wire[10:0] nl_Accum2_acc_1824_nl;
  wire[19:0] Product1_1_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_569_nl;
  wire[17:0] nl_Accum2_acc_569_nl;
  wire[15:0] Accum2_acc_563_nl;
  wire[16:0] nl_Accum2_acc_563_nl;
  wire[19:0] Product1_2_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_562_nl;
  wire[16:0] nl_Accum2_acc_562_nl;
  wire[19:0] Product1_4_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_561_nl;
  wire[16:0] nl_Accum2_acc_561_nl;
  wire[19:0] Product1_6_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_560_nl;
  wire[16:0] nl_Accum2_acc_560_nl;
  wire[19:0] Product1_8_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_568_nl;
  wire[16:0] nl_Accum2_acc_568_nl;
  wire[15:0] Accum2_acc_565_nl;
  wire[16:0] nl_Accum2_acc_565_nl;
  wire[15:0] Accum2_acc_559_nl;
  wire[16:0] nl_Accum2_acc_559_nl;
  wire[19:0] Product1_10_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_558_nl;
  wire[16:0] nl_Accum2_acc_558_nl;
  wire[19:0] Product1_12_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_564_nl;
  wire[16:0] nl_Accum2_acc_564_nl;
  wire[9:0] Accum2_acc_1825_nl;
  wire[10:0] nl_Accum2_acc_1825_nl;
  wire[19:0] Product1_1_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_582_nl;
  wire[17:0] nl_Accum2_acc_582_nl;
  wire[15:0] Accum2_acc_576_nl;
  wire[16:0] nl_Accum2_acc_576_nl;
  wire[19:0] Product1_2_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_575_nl;
  wire[16:0] nl_Accum2_acc_575_nl;
  wire[19:0] Product1_4_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_574_nl;
  wire[16:0] nl_Accum2_acc_574_nl;
  wire[19:0] Product1_6_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_573_nl;
  wire[16:0] nl_Accum2_acc_573_nl;
  wire[19:0] Product1_8_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_581_nl;
  wire[16:0] nl_Accum2_acc_581_nl;
  wire[15:0] Accum2_acc_578_nl;
  wire[16:0] nl_Accum2_acc_578_nl;
  wire[15:0] Accum2_acc_572_nl;
  wire[16:0] nl_Accum2_acc_572_nl;
  wire[19:0] Product1_10_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_571_nl;
  wire[16:0] nl_Accum2_acc_571_nl;
  wire[19:0] Product1_12_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_577_nl;
  wire[16:0] nl_Accum2_acc_577_nl;
  wire[9:0] Accum2_acc_1826_nl;
  wire[10:0] nl_Accum2_acc_1826_nl;
  wire[19:0] Product1_1_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_595_nl;
  wire[17:0] nl_Accum2_acc_595_nl;
  wire[15:0] Accum2_acc_589_nl;
  wire[16:0] nl_Accum2_acc_589_nl;
  wire[19:0] Product1_2_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_588_nl;
  wire[16:0] nl_Accum2_acc_588_nl;
  wire[19:0] Product1_4_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_587_nl;
  wire[16:0] nl_Accum2_acc_587_nl;
  wire[19:0] Product1_6_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_586_nl;
  wire[16:0] nl_Accum2_acc_586_nl;
  wire[19:0] Product1_8_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_594_nl;
  wire[16:0] nl_Accum2_acc_594_nl;
  wire[15:0] Accum2_acc_591_nl;
  wire[16:0] nl_Accum2_acc_591_nl;
  wire[15:0] Accum2_acc_585_nl;
  wire[16:0] nl_Accum2_acc_585_nl;
  wire[19:0] Product1_10_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_584_nl;
  wire[16:0] nl_Accum2_acc_584_nl;
  wire[19:0] Product1_12_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_590_nl;
  wire[16:0] nl_Accum2_acc_590_nl;
  wire[9:0] Accum2_acc_1827_nl;
  wire[10:0] nl_Accum2_acc_1827_nl;
  wire[19:0] Product1_1_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_608_nl;
  wire[17:0] nl_Accum2_acc_608_nl;
  wire[15:0] Accum2_acc_602_nl;
  wire[16:0] nl_Accum2_acc_602_nl;
  wire[19:0] Product1_2_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_601_nl;
  wire[16:0] nl_Accum2_acc_601_nl;
  wire[19:0] Product1_4_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_600_nl;
  wire[16:0] nl_Accum2_acc_600_nl;
  wire[19:0] Product1_6_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_599_nl;
  wire[16:0] nl_Accum2_acc_599_nl;
  wire[19:0] Product1_8_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_607_nl;
  wire[16:0] nl_Accum2_acc_607_nl;
  wire[15:0] Accum2_acc_604_nl;
  wire[16:0] nl_Accum2_acc_604_nl;
  wire[15:0] Accum2_acc_598_nl;
  wire[16:0] nl_Accum2_acc_598_nl;
  wire[19:0] Product1_10_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_597_nl;
  wire[16:0] nl_Accum2_acc_597_nl;
  wire[19:0] Product1_12_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_603_nl;
  wire[16:0] nl_Accum2_acc_603_nl;
  wire[9:0] Accum2_acc_1828_nl;
  wire[10:0] nl_Accum2_acc_1828_nl;
  wire[19:0] Product1_1_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_621_nl;
  wire[17:0] nl_Accum2_acc_621_nl;
  wire[15:0] Accum2_acc_615_nl;
  wire[16:0] nl_Accum2_acc_615_nl;
  wire[19:0] Product1_2_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_614_nl;
  wire[16:0] nl_Accum2_acc_614_nl;
  wire[19:0] Product1_4_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_613_nl;
  wire[16:0] nl_Accum2_acc_613_nl;
  wire[19:0] Product1_6_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_612_nl;
  wire[16:0] nl_Accum2_acc_612_nl;
  wire[19:0] Product1_8_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_620_nl;
  wire[16:0] nl_Accum2_acc_620_nl;
  wire[15:0] Accum2_acc_617_nl;
  wire[16:0] nl_Accum2_acc_617_nl;
  wire[15:0] Accum2_acc_611_nl;
  wire[16:0] nl_Accum2_acc_611_nl;
  wire[19:0] Product1_10_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_610_nl;
  wire[16:0] nl_Accum2_acc_610_nl;
  wire[19:0] Product1_12_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_616_nl;
  wire[16:0] nl_Accum2_acc_616_nl;
  wire[9:0] Accum2_acc_1829_nl;
  wire[10:0] nl_Accum2_acc_1829_nl;
  wire[19:0] Product1_1_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_634_nl;
  wire[17:0] nl_Accum2_acc_634_nl;
  wire[15:0] Accum2_acc_628_nl;
  wire[16:0] nl_Accum2_acc_628_nl;
  wire[19:0] Product1_2_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_627_nl;
  wire[16:0] nl_Accum2_acc_627_nl;
  wire[19:0] Product1_4_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_626_nl;
  wire[16:0] nl_Accum2_acc_626_nl;
  wire[19:0] Product1_6_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_625_nl;
  wire[16:0] nl_Accum2_acc_625_nl;
  wire[19:0] Product1_8_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_633_nl;
  wire[16:0] nl_Accum2_acc_633_nl;
  wire[15:0] Accum2_acc_630_nl;
  wire[16:0] nl_Accum2_acc_630_nl;
  wire[15:0] Accum2_acc_624_nl;
  wire[16:0] nl_Accum2_acc_624_nl;
  wire[19:0] Product1_10_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_623_nl;
  wire[16:0] nl_Accum2_acc_623_nl;
  wire[19:0] Product1_12_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_629_nl;
  wire[16:0] nl_Accum2_acc_629_nl;
  wire[9:0] Accum2_acc_1830_nl;
  wire[10:0] nl_Accum2_acc_1830_nl;
  wire[19:0] Product1_1_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_647_nl;
  wire[17:0] nl_Accum2_acc_647_nl;
  wire[15:0] Accum2_acc_641_nl;
  wire[16:0] nl_Accum2_acc_641_nl;
  wire[19:0] Product1_2_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_640_nl;
  wire[16:0] nl_Accum2_acc_640_nl;
  wire[19:0] Product1_4_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_639_nl;
  wire[16:0] nl_Accum2_acc_639_nl;
  wire[19:0] Product1_6_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_638_nl;
  wire[16:0] nl_Accum2_acc_638_nl;
  wire[19:0] Product1_8_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_646_nl;
  wire[16:0] nl_Accum2_acc_646_nl;
  wire[15:0] Accum2_acc_643_nl;
  wire[16:0] nl_Accum2_acc_643_nl;
  wire[15:0] Accum2_acc_637_nl;
  wire[16:0] nl_Accum2_acc_637_nl;
  wire[19:0] Product1_10_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_636_nl;
  wire[16:0] nl_Accum2_acc_636_nl;
  wire[19:0] Product1_12_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_642_nl;
  wire[16:0] nl_Accum2_acc_642_nl;
  wire[9:0] Accum2_acc_1831_nl;
  wire[10:0] nl_Accum2_acc_1831_nl;
  wire[19:0] Product1_1_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_660_nl;
  wire[17:0] nl_Accum2_acc_660_nl;
  wire[15:0] Accum2_acc_654_nl;
  wire[16:0] nl_Accum2_acc_654_nl;
  wire[19:0] Product1_2_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_653_nl;
  wire[16:0] nl_Accum2_acc_653_nl;
  wire[19:0] Product1_4_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_652_nl;
  wire[16:0] nl_Accum2_acc_652_nl;
  wire[19:0] Product1_6_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_651_nl;
  wire[16:0] nl_Accum2_acc_651_nl;
  wire[19:0] Product1_8_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_659_nl;
  wire[16:0] nl_Accum2_acc_659_nl;
  wire[15:0] Accum2_acc_656_nl;
  wire[16:0] nl_Accum2_acc_656_nl;
  wire[15:0] Accum2_acc_650_nl;
  wire[16:0] nl_Accum2_acc_650_nl;
  wire[19:0] Product1_10_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_649_nl;
  wire[16:0] nl_Accum2_acc_649_nl;
  wire[19:0] Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_655_nl;
  wire[16:0] nl_Accum2_acc_655_nl;
  wire[9:0] Accum2_acc_1832_nl;
  wire[10:0] nl_Accum2_acc_1832_nl;
  wire[19:0] Product1_1_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_673_nl;
  wire[17:0] nl_Accum2_acc_673_nl;
  wire[15:0] Accum2_acc_667_nl;
  wire[16:0] nl_Accum2_acc_667_nl;
  wire[19:0] Product1_2_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_666_nl;
  wire[16:0] nl_Accum2_acc_666_nl;
  wire[19:0] Product1_4_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_665_nl;
  wire[16:0] nl_Accum2_acc_665_nl;
  wire[19:0] Product1_6_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_664_nl;
  wire[16:0] nl_Accum2_acc_664_nl;
  wire[19:0] Product1_8_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_672_nl;
  wire[16:0] nl_Accum2_acc_672_nl;
  wire[15:0] Accum2_acc_669_nl;
  wire[16:0] nl_Accum2_acc_669_nl;
  wire[15:0] Accum2_acc_663_nl;
  wire[16:0] nl_Accum2_acc_663_nl;
  wire[19:0] Product1_10_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_662_nl;
  wire[16:0] nl_Accum2_acc_662_nl;
  wire[19:0] Product1_12_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_668_nl;
  wire[16:0] nl_Accum2_acc_668_nl;
  wire[9:0] Accum2_acc_1833_nl;
  wire[10:0] nl_Accum2_acc_1833_nl;
  wire[19:0] Product1_1_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_686_nl;
  wire[17:0] nl_Accum2_acc_686_nl;
  wire[15:0] Accum2_acc_680_nl;
  wire[16:0] nl_Accum2_acc_680_nl;
  wire[19:0] Product1_2_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_679_nl;
  wire[16:0] nl_Accum2_acc_679_nl;
  wire[19:0] Product1_4_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_678_nl;
  wire[16:0] nl_Accum2_acc_678_nl;
  wire[19:0] Product1_6_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_677_nl;
  wire[16:0] nl_Accum2_acc_677_nl;
  wire[19:0] Product1_8_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_685_nl;
  wire[16:0] nl_Accum2_acc_685_nl;
  wire[15:0] Accum2_acc_682_nl;
  wire[16:0] nl_Accum2_acc_682_nl;
  wire[15:0] Accum2_acc_676_nl;
  wire[16:0] nl_Accum2_acc_676_nl;
  wire[19:0] Product1_10_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_675_nl;
  wire[16:0] nl_Accum2_acc_675_nl;
  wire[19:0] Product1_12_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_681_nl;
  wire[16:0] nl_Accum2_acc_681_nl;
  wire[9:0] Accum2_acc_1834_nl;
  wire[10:0] nl_Accum2_acc_1834_nl;
  wire[19:0] Product1_1_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_699_nl;
  wire[17:0] nl_Accum2_acc_699_nl;
  wire[15:0] Accum2_acc_693_nl;
  wire[16:0] nl_Accum2_acc_693_nl;
  wire[19:0] Product1_2_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_692_nl;
  wire[16:0] nl_Accum2_acc_692_nl;
  wire[19:0] Product1_4_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_691_nl;
  wire[16:0] nl_Accum2_acc_691_nl;
  wire[19:0] Product1_6_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_690_nl;
  wire[16:0] nl_Accum2_acc_690_nl;
  wire[19:0] Product1_8_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_698_nl;
  wire[16:0] nl_Accum2_acc_698_nl;
  wire[15:0] Accum2_acc_695_nl;
  wire[16:0] nl_Accum2_acc_695_nl;
  wire[15:0] Accum2_acc_689_nl;
  wire[16:0] nl_Accum2_acc_689_nl;
  wire[19:0] Product1_10_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_688_nl;
  wire[16:0] nl_Accum2_acc_688_nl;
  wire[19:0] Product1_12_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_694_nl;
  wire[16:0] nl_Accum2_acc_694_nl;
  wire[9:0] Accum2_acc_1835_nl;
  wire[10:0] nl_Accum2_acc_1835_nl;
  wire[19:0] Product1_1_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_712_nl;
  wire[17:0] nl_Accum2_acc_712_nl;
  wire[15:0] Accum2_acc_706_nl;
  wire[16:0] nl_Accum2_acc_706_nl;
  wire[19:0] Product1_2_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_705_nl;
  wire[16:0] nl_Accum2_acc_705_nl;
  wire[19:0] Product1_4_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_704_nl;
  wire[16:0] nl_Accum2_acc_704_nl;
  wire[19:0] Product1_6_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_703_nl;
  wire[16:0] nl_Accum2_acc_703_nl;
  wire[19:0] Product1_8_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_711_nl;
  wire[16:0] nl_Accum2_acc_711_nl;
  wire[15:0] Accum2_acc_708_nl;
  wire[16:0] nl_Accum2_acc_708_nl;
  wire[15:0] Accum2_acc_702_nl;
  wire[16:0] nl_Accum2_acc_702_nl;
  wire[19:0] Product1_10_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_701_nl;
  wire[16:0] nl_Accum2_acc_701_nl;
  wire[19:0] Product1_12_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_707_nl;
  wire[16:0] nl_Accum2_acc_707_nl;
  wire[9:0] Accum2_acc_1836_nl;
  wire[10:0] nl_Accum2_acc_1836_nl;
  wire[19:0] Product1_1_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_725_nl;
  wire[17:0] nl_Accum2_acc_725_nl;
  wire[15:0] Accum2_acc_719_nl;
  wire[16:0] nl_Accum2_acc_719_nl;
  wire[19:0] Product1_2_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_718_nl;
  wire[16:0] nl_Accum2_acc_718_nl;
  wire[19:0] Product1_4_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_717_nl;
  wire[16:0] nl_Accum2_acc_717_nl;
  wire[19:0] Product1_6_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_716_nl;
  wire[16:0] nl_Accum2_acc_716_nl;
  wire[19:0] Product1_8_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_724_nl;
  wire[16:0] nl_Accum2_acc_724_nl;
  wire[15:0] Accum2_acc_721_nl;
  wire[16:0] nl_Accum2_acc_721_nl;
  wire[15:0] Accum2_acc_715_nl;
  wire[16:0] nl_Accum2_acc_715_nl;
  wire[19:0] Product1_10_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_714_nl;
  wire[16:0] nl_Accum2_acc_714_nl;
  wire[19:0] Product1_12_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_720_nl;
  wire[16:0] nl_Accum2_acc_720_nl;
  wire[9:0] Accum2_acc_1837_nl;
  wire[10:0] nl_Accum2_acc_1837_nl;
  wire[19:0] Product1_1_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_738_nl;
  wire[17:0] nl_Accum2_acc_738_nl;
  wire[15:0] Accum2_acc_732_nl;
  wire[16:0] nl_Accum2_acc_732_nl;
  wire[19:0] Product1_2_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_731_nl;
  wire[16:0] nl_Accum2_acc_731_nl;
  wire[19:0] Product1_4_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_730_nl;
  wire[16:0] nl_Accum2_acc_730_nl;
  wire[19:0] Product1_6_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_729_nl;
  wire[16:0] nl_Accum2_acc_729_nl;
  wire[19:0] Product1_8_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_737_nl;
  wire[16:0] nl_Accum2_acc_737_nl;
  wire[15:0] Accum2_acc_734_nl;
  wire[16:0] nl_Accum2_acc_734_nl;
  wire[15:0] Accum2_acc_728_nl;
  wire[16:0] nl_Accum2_acc_728_nl;
  wire[19:0] Product1_10_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_727_nl;
  wire[16:0] nl_Accum2_acc_727_nl;
  wire[19:0] Product1_12_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_733_nl;
  wire[16:0] nl_Accum2_acc_733_nl;
  wire[9:0] Accum2_acc_1838_nl;
  wire[10:0] nl_Accum2_acc_1838_nl;
  wire[19:0] Product1_1_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_751_nl;
  wire[17:0] nl_Accum2_acc_751_nl;
  wire[15:0] Accum2_acc_745_nl;
  wire[16:0] nl_Accum2_acc_745_nl;
  wire[19:0] Product1_2_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_744_nl;
  wire[16:0] nl_Accum2_acc_744_nl;
  wire[19:0] Product1_4_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_743_nl;
  wire[16:0] nl_Accum2_acc_743_nl;
  wire[19:0] Product1_6_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_742_nl;
  wire[16:0] nl_Accum2_acc_742_nl;
  wire[19:0] Product1_8_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_750_nl;
  wire[16:0] nl_Accum2_acc_750_nl;
  wire[15:0] Accum2_acc_747_nl;
  wire[16:0] nl_Accum2_acc_747_nl;
  wire[15:0] Accum2_acc_741_nl;
  wire[16:0] nl_Accum2_acc_741_nl;
  wire[19:0] Product1_10_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_740_nl;
  wire[16:0] nl_Accum2_acc_740_nl;
  wire[19:0] Product1_12_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_746_nl;
  wire[16:0] nl_Accum2_acc_746_nl;
  wire[9:0] Accum2_acc_1839_nl;
  wire[10:0] nl_Accum2_acc_1839_nl;
  wire[19:0] Product1_1_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_764_nl;
  wire[17:0] nl_Accum2_acc_764_nl;
  wire[15:0] Accum2_acc_758_nl;
  wire[16:0] nl_Accum2_acc_758_nl;
  wire[19:0] Product1_2_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_757_nl;
  wire[16:0] nl_Accum2_acc_757_nl;
  wire[19:0] Product1_4_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_756_nl;
  wire[16:0] nl_Accum2_acc_756_nl;
  wire[19:0] Product1_6_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_755_nl;
  wire[16:0] nl_Accum2_acc_755_nl;
  wire[19:0] Product1_8_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_763_nl;
  wire[16:0] nl_Accum2_acc_763_nl;
  wire[15:0] Accum2_acc_760_nl;
  wire[16:0] nl_Accum2_acc_760_nl;
  wire[15:0] Accum2_acc_754_nl;
  wire[16:0] nl_Accum2_acc_754_nl;
  wire[19:0] Product1_10_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_753_nl;
  wire[16:0] nl_Accum2_acc_753_nl;
  wire[19:0] Product1_12_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_759_nl;
  wire[16:0] nl_Accum2_acc_759_nl;
  wire[9:0] Accum2_acc_1840_nl;
  wire[10:0] nl_Accum2_acc_1840_nl;
  wire[19:0] Product1_1_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_777_nl;
  wire[17:0] nl_Accum2_acc_777_nl;
  wire[15:0] Accum2_acc_771_nl;
  wire[16:0] nl_Accum2_acc_771_nl;
  wire[19:0] Product1_2_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_770_nl;
  wire[16:0] nl_Accum2_acc_770_nl;
  wire[19:0] Product1_4_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_769_nl;
  wire[16:0] nl_Accum2_acc_769_nl;
  wire[19:0] Product1_6_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_768_nl;
  wire[16:0] nl_Accum2_acc_768_nl;
  wire[19:0] Product1_8_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_776_nl;
  wire[16:0] nl_Accum2_acc_776_nl;
  wire[15:0] Accum2_acc_773_nl;
  wire[16:0] nl_Accum2_acc_773_nl;
  wire[15:0] Accum2_acc_767_nl;
  wire[16:0] nl_Accum2_acc_767_nl;
  wire[19:0] Product1_10_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_766_nl;
  wire[16:0] nl_Accum2_acc_766_nl;
  wire[19:0] Product1_12_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_772_nl;
  wire[16:0] nl_Accum2_acc_772_nl;
  wire[9:0] Accum2_acc_1841_nl;
  wire[10:0] nl_Accum2_acc_1841_nl;
  wire[19:0] Product1_1_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_790_nl;
  wire[17:0] nl_Accum2_acc_790_nl;
  wire[15:0] Accum2_acc_784_nl;
  wire[16:0] nl_Accum2_acc_784_nl;
  wire[19:0] Product1_2_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_783_nl;
  wire[16:0] nl_Accum2_acc_783_nl;
  wire[19:0] Product1_4_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_782_nl;
  wire[16:0] nl_Accum2_acc_782_nl;
  wire[19:0] Product1_6_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_781_nl;
  wire[16:0] nl_Accum2_acc_781_nl;
  wire[19:0] Product1_8_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_789_nl;
  wire[16:0] nl_Accum2_acc_789_nl;
  wire[15:0] Accum2_acc_786_nl;
  wire[16:0] nl_Accum2_acc_786_nl;
  wire[15:0] Accum2_acc_780_nl;
  wire[16:0] nl_Accum2_acc_780_nl;
  wire[19:0] Product1_10_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_779_nl;
  wire[16:0] nl_Accum2_acc_779_nl;
  wire[19:0] Product1_12_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_785_nl;
  wire[16:0] nl_Accum2_acc_785_nl;
  wire[9:0] Accum2_acc_1842_nl;
  wire[10:0] nl_Accum2_acc_1842_nl;
  wire[19:0] Product1_1_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_803_nl;
  wire[17:0] nl_Accum2_acc_803_nl;
  wire[15:0] Accum2_acc_797_nl;
  wire[16:0] nl_Accum2_acc_797_nl;
  wire[19:0] Product1_2_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_796_nl;
  wire[16:0] nl_Accum2_acc_796_nl;
  wire[19:0] Product1_4_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_795_nl;
  wire[16:0] nl_Accum2_acc_795_nl;
  wire[19:0] Product1_6_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_794_nl;
  wire[16:0] nl_Accum2_acc_794_nl;
  wire[19:0] Product1_8_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_802_nl;
  wire[16:0] nl_Accum2_acc_802_nl;
  wire[15:0] Accum2_acc_799_nl;
  wire[16:0] nl_Accum2_acc_799_nl;
  wire[15:0] Accum2_acc_793_nl;
  wire[16:0] nl_Accum2_acc_793_nl;
  wire[19:0] Product1_10_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_792_nl;
  wire[16:0] nl_Accum2_acc_792_nl;
  wire[19:0] Product1_12_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_798_nl;
  wire[16:0] nl_Accum2_acc_798_nl;
  wire[9:0] Accum2_acc_1843_nl;
  wire[10:0] nl_Accum2_acc_1843_nl;
  wire[19:0] Product1_1_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_816_nl;
  wire[17:0] nl_Accum2_acc_816_nl;
  wire[15:0] Accum2_acc_810_nl;
  wire[16:0] nl_Accum2_acc_810_nl;
  wire[19:0] Product1_2_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_809_nl;
  wire[16:0] nl_Accum2_acc_809_nl;
  wire[19:0] Product1_4_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_808_nl;
  wire[16:0] nl_Accum2_acc_808_nl;
  wire[19:0] Product1_6_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_807_nl;
  wire[16:0] nl_Accum2_acc_807_nl;
  wire[19:0] Product1_8_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_815_nl;
  wire[16:0] nl_Accum2_acc_815_nl;
  wire[15:0] Accum2_acc_812_nl;
  wire[16:0] nl_Accum2_acc_812_nl;
  wire[15:0] Accum2_acc_806_nl;
  wire[16:0] nl_Accum2_acc_806_nl;
  wire[19:0] Product1_10_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_805_nl;
  wire[16:0] nl_Accum2_acc_805_nl;
  wire[19:0] Product1_12_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_811_nl;
  wire[16:0] nl_Accum2_acc_811_nl;
  wire[9:0] Accum2_acc_1844_nl;
  wire[10:0] nl_Accum2_acc_1844_nl;
  wire[19:0] Product1_1_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_829_nl;
  wire[17:0] nl_Accum2_acc_829_nl;
  wire[15:0] Accum2_acc_823_nl;
  wire[16:0] nl_Accum2_acc_823_nl;
  wire[19:0] Product1_2_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_822_nl;
  wire[16:0] nl_Accum2_acc_822_nl;
  wire[19:0] Product1_4_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_821_nl;
  wire[16:0] nl_Accum2_acc_821_nl;
  wire[19:0] Product1_6_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_820_nl;
  wire[16:0] nl_Accum2_acc_820_nl;
  wire[19:0] Product1_8_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_828_nl;
  wire[16:0] nl_Accum2_acc_828_nl;
  wire[15:0] Accum2_acc_825_nl;
  wire[16:0] nl_Accum2_acc_825_nl;
  wire[15:0] Accum2_acc_819_nl;
  wire[16:0] nl_Accum2_acc_819_nl;
  wire[19:0] Product1_10_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_818_nl;
  wire[16:0] nl_Accum2_acc_818_nl;
  wire[19:0] Product1_12_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_824_nl;
  wire[16:0] nl_Accum2_acc_824_nl;
  wire[9:0] Accum2_acc_1845_nl;
  wire[10:0] nl_Accum2_acc_1845_nl;
  wire[19:0] Product1_1_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_842_nl;
  wire[17:0] nl_Accum2_acc_842_nl;
  wire[15:0] Accum2_acc_836_nl;
  wire[16:0] nl_Accum2_acc_836_nl;
  wire[19:0] Product1_2_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_835_nl;
  wire[16:0] nl_Accum2_acc_835_nl;
  wire[19:0] Product1_4_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_834_nl;
  wire[16:0] nl_Accum2_acc_834_nl;
  wire[19:0] Product1_6_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_833_nl;
  wire[16:0] nl_Accum2_acc_833_nl;
  wire[19:0] Product1_8_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_841_nl;
  wire[16:0] nl_Accum2_acc_841_nl;
  wire[15:0] Accum2_acc_838_nl;
  wire[16:0] nl_Accum2_acc_838_nl;
  wire[15:0] Accum2_acc_832_nl;
  wire[16:0] nl_Accum2_acc_832_nl;
  wire[19:0] Product1_10_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_831_nl;
  wire[16:0] nl_Accum2_acc_831_nl;
  wire[19:0] Product1_12_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_837_nl;
  wire[16:0] nl_Accum2_acc_837_nl;
  wire[9:0] Accum2_acc_1846_nl;
  wire[10:0] nl_Accum2_acc_1846_nl;
  wire[19:0] Product1_1_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_855_nl;
  wire[17:0] nl_Accum2_acc_855_nl;
  wire[15:0] Accum2_acc_849_nl;
  wire[16:0] nl_Accum2_acc_849_nl;
  wire[19:0] Product1_2_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_848_nl;
  wire[16:0] nl_Accum2_acc_848_nl;
  wire[19:0] Product1_4_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_847_nl;
  wire[16:0] nl_Accum2_acc_847_nl;
  wire[19:0] Product1_6_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_846_nl;
  wire[16:0] nl_Accum2_acc_846_nl;
  wire[19:0] Product1_8_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_854_nl;
  wire[16:0] nl_Accum2_acc_854_nl;
  wire[15:0] Accum2_acc_851_nl;
  wire[16:0] nl_Accum2_acc_851_nl;
  wire[15:0] Accum2_acc_845_nl;
  wire[16:0] nl_Accum2_acc_845_nl;
  wire[19:0] Product1_10_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_844_nl;
  wire[16:0] nl_Accum2_acc_844_nl;
  wire[19:0] Product1_12_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_850_nl;
  wire[16:0] nl_Accum2_acc_850_nl;
  wire[9:0] Accum2_acc_1847_nl;
  wire[10:0] nl_Accum2_acc_1847_nl;
  wire[19:0] Product1_1_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_868_nl;
  wire[17:0] nl_Accum2_acc_868_nl;
  wire[15:0] Accum2_acc_862_nl;
  wire[16:0] nl_Accum2_acc_862_nl;
  wire[19:0] Product1_2_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_861_nl;
  wire[16:0] nl_Accum2_acc_861_nl;
  wire[19:0] Product1_4_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_860_nl;
  wire[16:0] nl_Accum2_acc_860_nl;
  wire[19:0] Product1_6_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_859_nl;
  wire[16:0] nl_Accum2_acc_859_nl;
  wire[19:0] Product1_8_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_867_nl;
  wire[16:0] nl_Accum2_acc_867_nl;
  wire[15:0] Accum2_acc_864_nl;
  wire[16:0] nl_Accum2_acc_864_nl;
  wire[15:0] Accum2_acc_858_nl;
  wire[16:0] nl_Accum2_acc_858_nl;
  wire[19:0] Product1_10_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_857_nl;
  wire[16:0] nl_Accum2_acc_857_nl;
  wire[19:0] Product1_12_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_863_nl;
  wire[16:0] nl_Accum2_acc_863_nl;
  wire[9:0] Accum2_acc_1848_nl;
  wire[10:0] nl_Accum2_acc_1848_nl;
  wire[19:0] Product1_1_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_881_nl;
  wire[17:0] nl_Accum2_acc_881_nl;
  wire[15:0] Accum2_acc_875_nl;
  wire[16:0] nl_Accum2_acc_875_nl;
  wire[19:0] Product1_2_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_874_nl;
  wire[16:0] nl_Accum2_acc_874_nl;
  wire[19:0] Product1_4_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_873_nl;
  wire[16:0] nl_Accum2_acc_873_nl;
  wire[19:0] Product1_6_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_872_nl;
  wire[16:0] nl_Accum2_acc_872_nl;
  wire[19:0] Product1_8_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_880_nl;
  wire[16:0] nl_Accum2_acc_880_nl;
  wire[15:0] Accum2_acc_877_nl;
  wire[16:0] nl_Accum2_acc_877_nl;
  wire[15:0] Accum2_acc_871_nl;
  wire[16:0] nl_Accum2_acc_871_nl;
  wire[19:0] Product1_10_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_870_nl;
  wire[16:0] nl_Accum2_acc_870_nl;
  wire[19:0] Product1_12_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_876_nl;
  wire[16:0] nl_Accum2_acc_876_nl;
  wire[9:0] Accum2_acc_1849_nl;
  wire[10:0] nl_Accum2_acc_1849_nl;
  wire[19:0] Product1_1_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_894_nl;
  wire[17:0] nl_Accum2_acc_894_nl;
  wire[15:0] Accum2_acc_888_nl;
  wire[16:0] nl_Accum2_acc_888_nl;
  wire[19:0] Product1_2_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_887_nl;
  wire[16:0] nl_Accum2_acc_887_nl;
  wire[19:0] Product1_4_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_886_nl;
  wire[16:0] nl_Accum2_acc_886_nl;
  wire[19:0] Product1_6_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_885_nl;
  wire[16:0] nl_Accum2_acc_885_nl;
  wire[19:0] Product1_8_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_893_nl;
  wire[16:0] nl_Accum2_acc_893_nl;
  wire[15:0] Accum2_acc_890_nl;
  wire[16:0] nl_Accum2_acc_890_nl;
  wire[15:0] Accum2_acc_884_nl;
  wire[16:0] nl_Accum2_acc_884_nl;
  wire[19:0] Product1_10_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_883_nl;
  wire[16:0] nl_Accum2_acc_883_nl;
  wire[19:0] Product1_12_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_889_nl;
  wire[16:0] nl_Accum2_acc_889_nl;
  wire[9:0] Accum2_acc_1850_nl;
  wire[10:0] nl_Accum2_acc_1850_nl;
  wire[19:0] Product1_1_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_907_nl;
  wire[17:0] nl_Accum2_acc_907_nl;
  wire[15:0] Accum2_acc_901_nl;
  wire[16:0] nl_Accum2_acc_901_nl;
  wire[19:0] Product1_2_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_900_nl;
  wire[16:0] nl_Accum2_acc_900_nl;
  wire[19:0] Product1_4_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_899_nl;
  wire[16:0] nl_Accum2_acc_899_nl;
  wire[19:0] Product1_6_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_898_nl;
  wire[16:0] nl_Accum2_acc_898_nl;
  wire[19:0] Product1_8_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_906_nl;
  wire[16:0] nl_Accum2_acc_906_nl;
  wire[15:0] Accum2_acc_903_nl;
  wire[16:0] nl_Accum2_acc_903_nl;
  wire[15:0] Accum2_acc_897_nl;
  wire[16:0] nl_Accum2_acc_897_nl;
  wire[19:0] Product1_10_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_896_nl;
  wire[16:0] nl_Accum2_acc_896_nl;
  wire[19:0] Product1_12_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_902_nl;
  wire[16:0] nl_Accum2_acc_902_nl;
  wire[9:0] Accum2_acc_1851_nl;
  wire[10:0] nl_Accum2_acc_1851_nl;
  wire[19:0] Product1_1_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_920_nl;
  wire[17:0] nl_Accum2_acc_920_nl;
  wire[15:0] Accum2_acc_914_nl;
  wire[16:0] nl_Accum2_acc_914_nl;
  wire[19:0] Product1_2_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_913_nl;
  wire[16:0] nl_Accum2_acc_913_nl;
  wire[19:0] Product1_4_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_912_nl;
  wire[16:0] nl_Accum2_acc_912_nl;
  wire[19:0] Product1_6_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_911_nl;
  wire[16:0] nl_Accum2_acc_911_nl;
  wire[19:0] Product1_8_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_919_nl;
  wire[16:0] nl_Accum2_acc_919_nl;
  wire[15:0] Accum2_acc_916_nl;
  wire[16:0] nl_Accum2_acc_916_nl;
  wire[15:0] Accum2_acc_910_nl;
  wire[16:0] nl_Accum2_acc_910_nl;
  wire[19:0] Product1_10_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_909_nl;
  wire[16:0] nl_Accum2_acc_909_nl;
  wire[19:0] Product1_12_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_915_nl;
  wire[16:0] nl_Accum2_acc_915_nl;
  wire[9:0] Accum2_acc_1852_nl;
  wire[10:0] nl_Accum2_acc_1852_nl;
  wire[19:0] Product1_1_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_933_nl;
  wire[17:0] nl_Accum2_acc_933_nl;
  wire[15:0] Accum2_acc_927_nl;
  wire[16:0] nl_Accum2_acc_927_nl;
  wire[19:0] Product1_2_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_926_nl;
  wire[16:0] nl_Accum2_acc_926_nl;
  wire[19:0] Product1_4_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_925_nl;
  wire[16:0] nl_Accum2_acc_925_nl;
  wire[19:0] Product1_6_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_924_nl;
  wire[16:0] nl_Accum2_acc_924_nl;
  wire[19:0] Product1_8_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_932_nl;
  wire[16:0] nl_Accum2_acc_932_nl;
  wire[15:0] Accum2_acc_929_nl;
  wire[16:0] nl_Accum2_acc_929_nl;
  wire[15:0] Accum2_acc_923_nl;
  wire[16:0] nl_Accum2_acc_923_nl;
  wire[19:0] Product1_10_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_922_nl;
  wire[16:0] nl_Accum2_acc_922_nl;
  wire[19:0] Product1_12_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_928_nl;
  wire[16:0] nl_Accum2_acc_928_nl;
  wire[9:0] Accum2_acc_1853_nl;
  wire[10:0] nl_Accum2_acc_1853_nl;
  wire[19:0] Product1_1_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_946_nl;
  wire[17:0] nl_Accum2_acc_946_nl;
  wire[15:0] Accum2_acc_940_nl;
  wire[16:0] nl_Accum2_acc_940_nl;
  wire[19:0] Product1_2_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_939_nl;
  wire[16:0] nl_Accum2_acc_939_nl;
  wire[19:0] Product1_4_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_938_nl;
  wire[16:0] nl_Accum2_acc_938_nl;
  wire[19:0] Product1_6_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_937_nl;
  wire[16:0] nl_Accum2_acc_937_nl;
  wire[19:0] Product1_8_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_945_nl;
  wire[16:0] nl_Accum2_acc_945_nl;
  wire[15:0] Accum2_acc_942_nl;
  wire[16:0] nl_Accum2_acc_942_nl;
  wire[15:0] Accum2_acc_936_nl;
  wire[16:0] nl_Accum2_acc_936_nl;
  wire[19:0] Product1_10_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_935_nl;
  wire[16:0] nl_Accum2_acc_935_nl;
  wire[19:0] Product1_12_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_941_nl;
  wire[16:0] nl_Accum2_acc_941_nl;
  wire[9:0] Accum2_acc_1854_nl;
  wire[10:0] nl_Accum2_acc_1854_nl;
  wire[19:0] Product1_1_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_959_nl;
  wire[17:0] nl_Accum2_acc_959_nl;
  wire[15:0] Accum2_acc_953_nl;
  wire[16:0] nl_Accum2_acc_953_nl;
  wire[19:0] Product1_2_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_952_nl;
  wire[16:0] nl_Accum2_acc_952_nl;
  wire[19:0] Product1_4_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_951_nl;
  wire[16:0] nl_Accum2_acc_951_nl;
  wire[19:0] Product1_6_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_950_nl;
  wire[16:0] nl_Accum2_acc_950_nl;
  wire[19:0] Product1_8_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_958_nl;
  wire[16:0] nl_Accum2_acc_958_nl;
  wire[15:0] Accum2_acc_955_nl;
  wire[16:0] nl_Accum2_acc_955_nl;
  wire[15:0] Accum2_acc_949_nl;
  wire[16:0] nl_Accum2_acc_949_nl;
  wire[19:0] Product1_10_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_948_nl;
  wire[16:0] nl_Accum2_acc_948_nl;
  wire[19:0] Product1_12_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_954_nl;
  wire[16:0] nl_Accum2_acc_954_nl;
  wire[9:0] Accum2_acc_1855_nl;
  wire[10:0] nl_Accum2_acc_1855_nl;
  wire[19:0] Product1_1_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_972_nl;
  wire[17:0] nl_Accum2_acc_972_nl;
  wire[15:0] Accum2_acc_966_nl;
  wire[16:0] nl_Accum2_acc_966_nl;
  wire[19:0] Product1_2_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_965_nl;
  wire[16:0] nl_Accum2_acc_965_nl;
  wire[19:0] Product1_4_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_964_nl;
  wire[16:0] nl_Accum2_acc_964_nl;
  wire[19:0] Product1_6_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_963_nl;
  wire[16:0] nl_Accum2_acc_963_nl;
  wire[19:0] Product1_8_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_971_nl;
  wire[16:0] nl_Accum2_acc_971_nl;
  wire[15:0] Accum2_acc_968_nl;
  wire[16:0] nl_Accum2_acc_968_nl;
  wire[15:0] Accum2_acc_962_nl;
  wire[16:0] nl_Accum2_acc_962_nl;
  wire[19:0] Product1_10_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_961_nl;
  wire[16:0] nl_Accum2_acc_961_nl;
  wire[19:0] Product1_12_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_967_nl;
  wire[16:0] nl_Accum2_acc_967_nl;
  wire[9:0] Accum2_acc_1856_nl;
  wire[10:0] nl_Accum2_acc_1856_nl;
  wire[19:0] Product1_1_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_985_nl;
  wire[17:0] nl_Accum2_acc_985_nl;
  wire[15:0] Accum2_acc_979_nl;
  wire[16:0] nl_Accum2_acc_979_nl;
  wire[19:0] Product1_2_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_978_nl;
  wire[16:0] nl_Accum2_acc_978_nl;
  wire[19:0] Product1_4_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_977_nl;
  wire[16:0] nl_Accum2_acc_977_nl;
  wire[19:0] Product1_6_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_976_nl;
  wire[16:0] nl_Accum2_acc_976_nl;
  wire[19:0] Product1_8_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_984_nl;
  wire[16:0] nl_Accum2_acc_984_nl;
  wire[15:0] Accum2_acc_981_nl;
  wire[16:0] nl_Accum2_acc_981_nl;
  wire[15:0] Accum2_acc_975_nl;
  wire[16:0] nl_Accum2_acc_975_nl;
  wire[19:0] Product1_10_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_974_nl;
  wire[16:0] nl_Accum2_acc_974_nl;
  wire[19:0] Product1_12_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_980_nl;
  wire[16:0] nl_Accum2_acc_980_nl;
  wire[9:0] Accum2_acc_1857_nl;
  wire[10:0] nl_Accum2_acc_1857_nl;
  wire[19:0] Product1_1_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_998_nl;
  wire[17:0] nl_Accum2_acc_998_nl;
  wire[15:0] Accum2_acc_992_nl;
  wire[16:0] nl_Accum2_acc_992_nl;
  wire[19:0] Product1_2_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_991_nl;
  wire[16:0] nl_Accum2_acc_991_nl;
  wire[19:0] Product1_4_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_990_nl;
  wire[16:0] nl_Accum2_acc_990_nl;
  wire[19:0] Product1_6_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_989_nl;
  wire[16:0] nl_Accum2_acc_989_nl;
  wire[19:0] Product1_8_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_997_nl;
  wire[16:0] nl_Accum2_acc_997_nl;
  wire[15:0] Accum2_acc_994_nl;
  wire[16:0] nl_Accum2_acc_994_nl;
  wire[15:0] Accum2_acc_988_nl;
  wire[16:0] nl_Accum2_acc_988_nl;
  wire[19:0] Product1_10_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_987_nl;
  wire[16:0] nl_Accum2_acc_987_nl;
  wire[19:0] Product1_12_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_993_nl;
  wire[16:0] nl_Accum2_acc_993_nl;
  wire[9:0] Accum2_acc_1858_nl;
  wire[10:0] nl_Accum2_acc_1858_nl;
  wire[19:0] Product1_1_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1011_nl;
  wire[17:0] nl_Accum2_acc_1011_nl;
  wire[15:0] Accum2_acc_1005_nl;
  wire[16:0] nl_Accum2_acc_1005_nl;
  wire[19:0] Product1_2_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1004_nl;
  wire[16:0] nl_Accum2_acc_1004_nl;
  wire[19:0] Product1_4_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1003_nl;
  wire[16:0] nl_Accum2_acc_1003_nl;
  wire[19:0] Product1_6_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1002_nl;
  wire[16:0] nl_Accum2_acc_1002_nl;
  wire[19:0] Product1_8_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1010_nl;
  wire[16:0] nl_Accum2_acc_1010_nl;
  wire[15:0] Accum2_acc_1007_nl;
  wire[16:0] nl_Accum2_acc_1007_nl;
  wire[15:0] Accum2_acc_1001_nl;
  wire[16:0] nl_Accum2_acc_1001_nl;
  wire[19:0] Product1_10_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1000_nl;
  wire[16:0] nl_Accum2_acc_1000_nl;
  wire[19:0] Product1_12_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1006_nl;
  wire[16:0] nl_Accum2_acc_1006_nl;
  wire[9:0] Accum2_acc_1859_nl;
  wire[10:0] nl_Accum2_acc_1859_nl;
  wire[19:0] Product1_1_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1024_nl;
  wire[17:0] nl_Accum2_acc_1024_nl;
  wire[15:0] Accum2_acc_1018_nl;
  wire[16:0] nl_Accum2_acc_1018_nl;
  wire[19:0] Product1_2_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1017_nl;
  wire[16:0] nl_Accum2_acc_1017_nl;
  wire[19:0] Product1_4_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1016_nl;
  wire[16:0] nl_Accum2_acc_1016_nl;
  wire[19:0] Product1_6_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1015_nl;
  wire[16:0] nl_Accum2_acc_1015_nl;
  wire[19:0] Product1_8_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1023_nl;
  wire[16:0] nl_Accum2_acc_1023_nl;
  wire[15:0] Accum2_acc_1020_nl;
  wire[16:0] nl_Accum2_acc_1020_nl;
  wire[15:0] Accum2_acc_1014_nl;
  wire[16:0] nl_Accum2_acc_1014_nl;
  wire[19:0] Product1_10_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1013_nl;
  wire[16:0] nl_Accum2_acc_1013_nl;
  wire[19:0] Product1_12_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1019_nl;
  wire[16:0] nl_Accum2_acc_1019_nl;
  wire[9:0] Accum2_acc_1860_nl;
  wire[10:0] nl_Accum2_acc_1860_nl;
  wire[19:0] Product1_1_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1037_nl;
  wire[17:0] nl_Accum2_acc_1037_nl;
  wire[15:0] Accum2_acc_1031_nl;
  wire[16:0] nl_Accum2_acc_1031_nl;
  wire[19:0] Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1030_nl;
  wire[16:0] nl_Accum2_acc_1030_nl;
  wire[19:0] Product1_4_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1029_nl;
  wire[16:0] nl_Accum2_acc_1029_nl;
  wire[19:0] Product1_6_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1028_nl;
  wire[16:0] nl_Accum2_acc_1028_nl;
  wire[19:0] Product1_8_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1036_nl;
  wire[16:0] nl_Accum2_acc_1036_nl;
  wire[15:0] Accum2_acc_1033_nl;
  wire[16:0] nl_Accum2_acc_1033_nl;
  wire[15:0] Accum2_acc_1027_nl;
  wire[16:0] nl_Accum2_acc_1027_nl;
  wire[19:0] Product1_10_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1026_nl;
  wire[16:0] nl_Accum2_acc_1026_nl;
  wire[19:0] Product1_12_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1032_nl;
  wire[16:0] nl_Accum2_acc_1032_nl;
  wire[9:0] Accum2_acc_1861_nl;
  wire[10:0] nl_Accum2_acc_1861_nl;
  wire[19:0] Product1_1_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1050_nl;
  wire[17:0] nl_Accum2_acc_1050_nl;
  wire[15:0] Accum2_acc_1044_nl;
  wire[16:0] nl_Accum2_acc_1044_nl;
  wire[19:0] Product1_2_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1043_nl;
  wire[16:0] nl_Accum2_acc_1043_nl;
  wire[19:0] Product1_4_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1042_nl;
  wire[16:0] nl_Accum2_acc_1042_nl;
  wire[19:0] Product1_6_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1041_nl;
  wire[16:0] nl_Accum2_acc_1041_nl;
  wire[19:0] Product1_8_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1049_nl;
  wire[16:0] nl_Accum2_acc_1049_nl;
  wire[15:0] Accum2_acc_1046_nl;
  wire[16:0] nl_Accum2_acc_1046_nl;
  wire[15:0] Accum2_acc_1040_nl;
  wire[16:0] nl_Accum2_acc_1040_nl;
  wire[19:0] Product1_10_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1039_nl;
  wire[16:0] nl_Accum2_acc_1039_nl;
  wire[19:0] Product1_12_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1045_nl;
  wire[16:0] nl_Accum2_acc_1045_nl;
  wire[9:0] Accum2_acc_1862_nl;
  wire[10:0] nl_Accum2_acc_1862_nl;
  wire[19:0] Product1_1_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1063_nl;
  wire[17:0] nl_Accum2_acc_1063_nl;
  wire[15:0] Accum2_acc_1057_nl;
  wire[16:0] nl_Accum2_acc_1057_nl;
  wire[19:0] Product1_2_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1056_nl;
  wire[16:0] nl_Accum2_acc_1056_nl;
  wire[19:0] Product1_4_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1055_nl;
  wire[16:0] nl_Accum2_acc_1055_nl;
  wire[19:0] Product1_6_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1054_nl;
  wire[16:0] nl_Accum2_acc_1054_nl;
  wire[19:0] Product1_8_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1062_nl;
  wire[16:0] nl_Accum2_acc_1062_nl;
  wire[15:0] Accum2_acc_1059_nl;
  wire[16:0] nl_Accum2_acc_1059_nl;
  wire[15:0] Accum2_acc_1053_nl;
  wire[16:0] nl_Accum2_acc_1053_nl;
  wire[19:0] Product1_10_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1052_nl;
  wire[16:0] nl_Accum2_acc_1052_nl;
  wire[19:0] Product1_12_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1058_nl;
  wire[16:0] nl_Accum2_acc_1058_nl;
  wire[9:0] Accum2_acc_1863_nl;
  wire[10:0] nl_Accum2_acc_1863_nl;
  wire[19:0] Product1_1_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1076_nl;
  wire[17:0] nl_Accum2_acc_1076_nl;
  wire[15:0] Accum2_acc_1070_nl;
  wire[16:0] nl_Accum2_acc_1070_nl;
  wire[19:0] Product1_2_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1069_nl;
  wire[16:0] nl_Accum2_acc_1069_nl;
  wire[19:0] Product1_4_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1068_nl;
  wire[16:0] nl_Accum2_acc_1068_nl;
  wire[19:0] Product1_6_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1067_nl;
  wire[16:0] nl_Accum2_acc_1067_nl;
  wire[19:0] Product1_8_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1075_nl;
  wire[16:0] nl_Accum2_acc_1075_nl;
  wire[15:0] Accum2_acc_1072_nl;
  wire[16:0] nl_Accum2_acc_1072_nl;
  wire[15:0] Accum2_acc_1066_nl;
  wire[16:0] nl_Accum2_acc_1066_nl;
  wire[19:0] Product1_10_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1065_nl;
  wire[16:0] nl_Accum2_acc_1065_nl;
  wire[19:0] Product1_12_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1071_nl;
  wire[16:0] nl_Accum2_acc_1071_nl;
  wire[9:0] Accum2_acc_1864_nl;
  wire[10:0] nl_Accum2_acc_1864_nl;
  wire[19:0] Product1_1_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1089_nl;
  wire[17:0] nl_Accum2_acc_1089_nl;
  wire[15:0] Accum2_acc_1083_nl;
  wire[16:0] nl_Accum2_acc_1083_nl;
  wire[19:0] Product1_2_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1082_nl;
  wire[16:0] nl_Accum2_acc_1082_nl;
  wire[19:0] Product1_4_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1081_nl;
  wire[16:0] nl_Accum2_acc_1081_nl;
  wire[19:0] Product1_6_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1080_nl;
  wire[16:0] nl_Accum2_acc_1080_nl;
  wire[19:0] Product1_8_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1088_nl;
  wire[16:0] nl_Accum2_acc_1088_nl;
  wire[15:0] Accum2_acc_1085_nl;
  wire[16:0] nl_Accum2_acc_1085_nl;
  wire[15:0] Accum2_acc_1079_nl;
  wire[16:0] nl_Accum2_acc_1079_nl;
  wire[19:0] Product1_10_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1078_nl;
  wire[16:0] nl_Accum2_acc_1078_nl;
  wire[19:0] Product1_12_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1084_nl;
  wire[16:0] nl_Accum2_acc_1084_nl;
  wire[9:0] Accum2_acc_1865_nl;
  wire[10:0] nl_Accum2_acc_1865_nl;
  wire[19:0] Product1_1_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1102_nl;
  wire[17:0] nl_Accum2_acc_1102_nl;
  wire[15:0] Accum2_acc_1096_nl;
  wire[16:0] nl_Accum2_acc_1096_nl;
  wire[19:0] Product1_2_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1095_nl;
  wire[16:0] nl_Accum2_acc_1095_nl;
  wire[19:0] Product1_4_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1094_nl;
  wire[16:0] nl_Accum2_acc_1094_nl;
  wire[19:0] Product1_6_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1093_nl;
  wire[16:0] nl_Accum2_acc_1093_nl;
  wire[19:0] Product1_8_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1101_nl;
  wire[16:0] nl_Accum2_acc_1101_nl;
  wire[15:0] Accum2_acc_1098_nl;
  wire[16:0] nl_Accum2_acc_1098_nl;
  wire[15:0] Accum2_acc_1092_nl;
  wire[16:0] nl_Accum2_acc_1092_nl;
  wire[19:0] Product1_10_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1091_nl;
  wire[16:0] nl_Accum2_acc_1091_nl;
  wire[19:0] Product1_12_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1097_nl;
  wire[16:0] nl_Accum2_acc_1097_nl;
  wire[9:0] Accum2_acc_1866_nl;
  wire[10:0] nl_Accum2_acc_1866_nl;
  wire[19:0] Product1_1_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1115_nl;
  wire[17:0] nl_Accum2_acc_1115_nl;
  wire[15:0] Accum2_acc_1109_nl;
  wire[16:0] nl_Accum2_acc_1109_nl;
  wire[19:0] Product1_2_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1108_nl;
  wire[16:0] nl_Accum2_acc_1108_nl;
  wire[19:0] Product1_4_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1107_nl;
  wire[16:0] nl_Accum2_acc_1107_nl;
  wire[19:0] Product1_6_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1106_nl;
  wire[16:0] nl_Accum2_acc_1106_nl;
  wire[19:0] Product1_8_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1114_nl;
  wire[16:0] nl_Accum2_acc_1114_nl;
  wire[15:0] Accum2_acc_1111_nl;
  wire[16:0] nl_Accum2_acc_1111_nl;
  wire[15:0] Accum2_acc_1105_nl;
  wire[16:0] nl_Accum2_acc_1105_nl;
  wire[19:0] Product1_10_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1104_nl;
  wire[16:0] nl_Accum2_acc_1104_nl;
  wire[19:0] Product1_12_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1110_nl;
  wire[16:0] nl_Accum2_acc_1110_nl;
  wire[9:0] Accum2_acc_1867_nl;
  wire[10:0] nl_Accum2_acc_1867_nl;
  wire[19:0] Product1_1_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1128_nl;
  wire[17:0] nl_Accum2_acc_1128_nl;
  wire[15:0] Accum2_acc_1122_nl;
  wire[16:0] nl_Accum2_acc_1122_nl;
  wire[19:0] Product1_2_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1121_nl;
  wire[16:0] nl_Accum2_acc_1121_nl;
  wire[19:0] Product1_4_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1120_nl;
  wire[16:0] nl_Accum2_acc_1120_nl;
  wire[19:0] Product1_6_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1119_nl;
  wire[16:0] nl_Accum2_acc_1119_nl;
  wire[19:0] Product1_8_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1127_nl;
  wire[16:0] nl_Accum2_acc_1127_nl;
  wire[15:0] Accum2_acc_1124_nl;
  wire[16:0] nl_Accum2_acc_1124_nl;
  wire[15:0] Accum2_acc_1118_nl;
  wire[16:0] nl_Accum2_acc_1118_nl;
  wire[19:0] Product1_10_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1117_nl;
  wire[16:0] nl_Accum2_acc_1117_nl;
  wire[19:0] Product1_12_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1123_nl;
  wire[16:0] nl_Accum2_acc_1123_nl;
  wire[9:0] Accum2_acc_1868_nl;
  wire[10:0] nl_Accum2_acc_1868_nl;
  wire[19:0] Product1_1_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1141_nl;
  wire[17:0] nl_Accum2_acc_1141_nl;
  wire[15:0] Accum2_acc_1135_nl;
  wire[16:0] nl_Accum2_acc_1135_nl;
  wire[19:0] Product1_2_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1134_nl;
  wire[16:0] nl_Accum2_acc_1134_nl;
  wire[19:0] Product1_4_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1133_nl;
  wire[16:0] nl_Accum2_acc_1133_nl;
  wire[19:0] Product1_6_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1132_nl;
  wire[16:0] nl_Accum2_acc_1132_nl;
  wire[19:0] Product1_8_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1140_nl;
  wire[16:0] nl_Accum2_acc_1140_nl;
  wire[15:0] Accum2_acc_1137_nl;
  wire[16:0] nl_Accum2_acc_1137_nl;
  wire[15:0] Accum2_acc_1131_nl;
  wire[16:0] nl_Accum2_acc_1131_nl;
  wire[19:0] Product1_10_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1130_nl;
  wire[16:0] nl_Accum2_acc_1130_nl;
  wire[19:0] Product1_12_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1136_nl;
  wire[16:0] nl_Accum2_acc_1136_nl;
  wire[9:0] Accum2_acc_1869_nl;
  wire[10:0] nl_Accum2_acc_1869_nl;
  wire[19:0] Product1_1_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1154_nl;
  wire[17:0] nl_Accum2_acc_1154_nl;
  wire[15:0] Accum2_acc_1148_nl;
  wire[16:0] nl_Accum2_acc_1148_nl;
  wire[19:0] Product1_2_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1147_nl;
  wire[16:0] nl_Accum2_acc_1147_nl;
  wire[19:0] Product1_4_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1146_nl;
  wire[16:0] nl_Accum2_acc_1146_nl;
  wire[19:0] Product1_6_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1145_nl;
  wire[16:0] nl_Accum2_acc_1145_nl;
  wire[19:0] Product1_8_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1153_nl;
  wire[16:0] nl_Accum2_acc_1153_nl;
  wire[15:0] Accum2_acc_1150_nl;
  wire[16:0] nl_Accum2_acc_1150_nl;
  wire[15:0] Accum2_acc_1144_nl;
  wire[16:0] nl_Accum2_acc_1144_nl;
  wire[19:0] Product1_10_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1143_nl;
  wire[16:0] nl_Accum2_acc_1143_nl;
  wire[19:0] Product1_12_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1149_nl;
  wire[16:0] nl_Accum2_acc_1149_nl;
  wire[9:0] Accum2_acc_1870_nl;
  wire[10:0] nl_Accum2_acc_1870_nl;
  wire[19:0] Product1_1_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1167_nl;
  wire[17:0] nl_Accum2_acc_1167_nl;
  wire[15:0] Accum2_acc_1161_nl;
  wire[16:0] nl_Accum2_acc_1161_nl;
  wire[19:0] Product1_2_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1160_nl;
  wire[16:0] nl_Accum2_acc_1160_nl;
  wire[19:0] Product1_4_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1159_nl;
  wire[16:0] nl_Accum2_acc_1159_nl;
  wire[19:0] Product1_6_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1158_nl;
  wire[16:0] nl_Accum2_acc_1158_nl;
  wire[19:0] Product1_8_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1166_nl;
  wire[16:0] nl_Accum2_acc_1166_nl;
  wire[15:0] Accum2_acc_1163_nl;
  wire[16:0] nl_Accum2_acc_1163_nl;
  wire[15:0] Accum2_acc_1157_nl;
  wire[16:0] nl_Accum2_acc_1157_nl;
  wire[19:0] Product1_10_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1156_nl;
  wire[16:0] nl_Accum2_acc_1156_nl;
  wire[19:0] Product1_12_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1162_nl;
  wire[16:0] nl_Accum2_acc_1162_nl;
  wire[9:0] Accum2_acc_1871_nl;
  wire[10:0] nl_Accum2_acc_1871_nl;
  wire[19:0] Product1_1_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1180_nl;
  wire[17:0] nl_Accum2_acc_1180_nl;
  wire[15:0] Accum2_acc_1174_nl;
  wire[16:0] nl_Accum2_acc_1174_nl;
  wire[19:0] Product1_2_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1173_nl;
  wire[16:0] nl_Accum2_acc_1173_nl;
  wire[19:0] Product1_4_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1172_nl;
  wire[16:0] nl_Accum2_acc_1172_nl;
  wire[19:0] Product1_6_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1171_nl;
  wire[16:0] nl_Accum2_acc_1171_nl;
  wire[19:0] Product1_8_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1179_nl;
  wire[16:0] nl_Accum2_acc_1179_nl;
  wire[15:0] Accum2_acc_1176_nl;
  wire[16:0] nl_Accum2_acc_1176_nl;
  wire[15:0] Accum2_acc_1170_nl;
  wire[16:0] nl_Accum2_acc_1170_nl;
  wire[19:0] Product1_10_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1169_nl;
  wire[16:0] nl_Accum2_acc_1169_nl;
  wire[19:0] Product1_12_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1175_nl;
  wire[16:0] nl_Accum2_acc_1175_nl;
  wire[9:0] Accum2_acc_1872_nl;
  wire[10:0] nl_Accum2_acc_1872_nl;
  wire[19:0] Product1_1_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1193_nl;
  wire[17:0] nl_Accum2_acc_1193_nl;
  wire[15:0] Accum2_acc_1187_nl;
  wire[16:0] nl_Accum2_acc_1187_nl;
  wire[19:0] Product1_2_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1186_nl;
  wire[16:0] nl_Accum2_acc_1186_nl;
  wire[19:0] Product1_4_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1185_nl;
  wire[16:0] nl_Accum2_acc_1185_nl;
  wire[19:0] Product1_6_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1184_nl;
  wire[16:0] nl_Accum2_acc_1184_nl;
  wire[19:0] Product1_8_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1192_nl;
  wire[16:0] nl_Accum2_acc_1192_nl;
  wire[15:0] Accum2_acc_1189_nl;
  wire[16:0] nl_Accum2_acc_1189_nl;
  wire[15:0] Accum2_acc_1183_nl;
  wire[16:0] nl_Accum2_acc_1183_nl;
  wire[19:0] Product1_10_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1182_nl;
  wire[16:0] nl_Accum2_acc_1182_nl;
  wire[19:0] Product1_12_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1188_nl;
  wire[16:0] nl_Accum2_acc_1188_nl;
  wire[9:0] Accum2_acc_1873_nl;
  wire[10:0] nl_Accum2_acc_1873_nl;
  wire[19:0] Product1_1_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1206_nl;
  wire[17:0] nl_Accum2_acc_1206_nl;
  wire[15:0] Accum2_acc_1200_nl;
  wire[16:0] nl_Accum2_acc_1200_nl;
  wire[19:0] Product1_2_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1199_nl;
  wire[16:0] nl_Accum2_acc_1199_nl;
  wire[19:0] Product1_4_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1198_nl;
  wire[16:0] nl_Accum2_acc_1198_nl;
  wire[19:0] Product1_6_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1197_nl;
  wire[16:0] nl_Accum2_acc_1197_nl;
  wire[19:0] Product1_8_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1205_nl;
  wire[16:0] nl_Accum2_acc_1205_nl;
  wire[15:0] Accum2_acc_1202_nl;
  wire[16:0] nl_Accum2_acc_1202_nl;
  wire[15:0] Accum2_acc_1196_nl;
  wire[16:0] nl_Accum2_acc_1196_nl;
  wire[19:0] Product1_10_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1195_nl;
  wire[16:0] nl_Accum2_acc_1195_nl;
  wire[19:0] Product1_12_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1201_nl;
  wire[16:0] nl_Accum2_acc_1201_nl;
  wire[9:0] Accum2_acc_1874_nl;
  wire[10:0] nl_Accum2_acc_1874_nl;
  wire[19:0] Product1_1_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1219_nl;
  wire[17:0] nl_Accum2_acc_1219_nl;
  wire[15:0] Accum2_acc_1213_nl;
  wire[16:0] nl_Accum2_acc_1213_nl;
  wire[19:0] Product1_2_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1212_nl;
  wire[16:0] nl_Accum2_acc_1212_nl;
  wire[19:0] Product1_4_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1211_nl;
  wire[16:0] nl_Accum2_acc_1211_nl;
  wire[19:0] Product1_6_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1210_nl;
  wire[16:0] nl_Accum2_acc_1210_nl;
  wire[19:0] Product1_8_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1218_nl;
  wire[16:0] nl_Accum2_acc_1218_nl;
  wire[15:0] Accum2_acc_1215_nl;
  wire[16:0] nl_Accum2_acc_1215_nl;
  wire[15:0] Accum2_acc_1209_nl;
  wire[16:0] nl_Accum2_acc_1209_nl;
  wire[19:0] Product1_10_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1208_nl;
  wire[16:0] nl_Accum2_acc_1208_nl;
  wire[19:0] Product1_12_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1214_nl;
  wire[16:0] nl_Accum2_acc_1214_nl;
  wire[9:0] Accum2_acc_1875_nl;
  wire[10:0] nl_Accum2_acc_1875_nl;
  wire[19:0] Product1_1_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1232_nl;
  wire[17:0] nl_Accum2_acc_1232_nl;
  wire[15:0] Accum2_acc_1226_nl;
  wire[16:0] nl_Accum2_acc_1226_nl;
  wire[19:0] Product1_2_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1225_nl;
  wire[16:0] nl_Accum2_acc_1225_nl;
  wire[19:0] Product1_4_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1224_nl;
  wire[16:0] nl_Accum2_acc_1224_nl;
  wire[19:0] Product1_6_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1223_nl;
  wire[16:0] nl_Accum2_acc_1223_nl;
  wire[19:0] Product1_8_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1231_nl;
  wire[16:0] nl_Accum2_acc_1231_nl;
  wire[15:0] Accum2_acc_1228_nl;
  wire[16:0] nl_Accum2_acc_1228_nl;
  wire[15:0] Accum2_acc_1222_nl;
  wire[16:0] nl_Accum2_acc_1222_nl;
  wire[19:0] Product1_10_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1221_nl;
  wire[16:0] nl_Accum2_acc_1221_nl;
  wire[19:0] Product1_12_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1227_nl;
  wire[16:0] nl_Accum2_acc_1227_nl;
  wire[9:0] Accum2_acc_1876_nl;
  wire[10:0] nl_Accum2_acc_1876_nl;
  wire[19:0] Product1_1_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1245_nl;
  wire[17:0] nl_Accum2_acc_1245_nl;
  wire[15:0] Accum2_acc_1239_nl;
  wire[16:0] nl_Accum2_acc_1239_nl;
  wire[19:0] Product1_2_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1238_nl;
  wire[16:0] nl_Accum2_acc_1238_nl;
  wire[19:0] Product1_4_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1237_nl;
  wire[16:0] nl_Accum2_acc_1237_nl;
  wire[19:0] Product1_6_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1236_nl;
  wire[16:0] nl_Accum2_acc_1236_nl;
  wire[19:0] Product1_8_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1244_nl;
  wire[16:0] nl_Accum2_acc_1244_nl;
  wire[15:0] Accum2_acc_1241_nl;
  wire[16:0] nl_Accum2_acc_1241_nl;
  wire[15:0] Accum2_acc_1235_nl;
  wire[16:0] nl_Accum2_acc_1235_nl;
  wire[19:0] Product1_10_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1234_nl;
  wire[16:0] nl_Accum2_acc_1234_nl;
  wire[19:0] Product1_12_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1240_nl;
  wire[16:0] nl_Accum2_acc_1240_nl;
  wire[9:0] Accum2_acc_1877_nl;
  wire[10:0] nl_Accum2_acc_1877_nl;
  wire[19:0] Product1_1_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1258_nl;
  wire[17:0] nl_Accum2_acc_1258_nl;
  wire[15:0] Accum2_acc_1252_nl;
  wire[16:0] nl_Accum2_acc_1252_nl;
  wire[19:0] Product1_2_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1251_nl;
  wire[16:0] nl_Accum2_acc_1251_nl;
  wire[19:0] Product1_4_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1250_nl;
  wire[16:0] nl_Accum2_acc_1250_nl;
  wire[19:0] Product1_6_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1249_nl;
  wire[16:0] nl_Accum2_acc_1249_nl;
  wire[19:0] Product1_8_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1257_nl;
  wire[16:0] nl_Accum2_acc_1257_nl;
  wire[15:0] Accum2_acc_1254_nl;
  wire[16:0] nl_Accum2_acc_1254_nl;
  wire[15:0] Accum2_acc_1248_nl;
  wire[16:0] nl_Accum2_acc_1248_nl;
  wire[19:0] Product1_10_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1247_nl;
  wire[16:0] nl_Accum2_acc_1247_nl;
  wire[19:0] Product1_12_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1253_nl;
  wire[16:0] nl_Accum2_acc_1253_nl;
  wire[9:0] Accum2_acc_1878_nl;
  wire[10:0] nl_Accum2_acc_1878_nl;
  wire[19:0] Product1_1_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1271_nl;
  wire[17:0] nl_Accum2_acc_1271_nl;
  wire[15:0] Accum2_acc_1265_nl;
  wire[16:0] nl_Accum2_acc_1265_nl;
  wire[19:0] Product1_2_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1264_nl;
  wire[16:0] nl_Accum2_acc_1264_nl;
  wire[19:0] Product1_4_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1263_nl;
  wire[16:0] nl_Accum2_acc_1263_nl;
  wire[19:0] Product1_6_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1262_nl;
  wire[16:0] nl_Accum2_acc_1262_nl;
  wire[19:0] Product1_8_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1270_nl;
  wire[16:0] nl_Accum2_acc_1270_nl;
  wire[15:0] Accum2_acc_1267_nl;
  wire[16:0] nl_Accum2_acc_1267_nl;
  wire[15:0] Accum2_acc_1261_nl;
  wire[16:0] nl_Accum2_acc_1261_nl;
  wire[19:0] Product1_10_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1260_nl;
  wire[16:0] nl_Accum2_acc_1260_nl;
  wire[19:0] Product1_12_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1266_nl;
  wire[16:0] nl_Accum2_acc_1266_nl;
  wire[9:0] Accum2_acc_1879_nl;
  wire[10:0] nl_Accum2_acc_1879_nl;
  wire[19:0] Product1_1_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1284_nl;
  wire[17:0] nl_Accum2_acc_1284_nl;
  wire[15:0] Accum2_acc_1278_nl;
  wire[16:0] nl_Accum2_acc_1278_nl;
  wire[19:0] Product1_2_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1277_nl;
  wire[16:0] nl_Accum2_acc_1277_nl;
  wire[19:0] Product1_4_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1276_nl;
  wire[16:0] nl_Accum2_acc_1276_nl;
  wire[19:0] Product1_6_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1275_nl;
  wire[16:0] nl_Accum2_acc_1275_nl;
  wire[19:0] Product1_8_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1283_nl;
  wire[16:0] nl_Accum2_acc_1283_nl;
  wire[15:0] Accum2_acc_1280_nl;
  wire[16:0] nl_Accum2_acc_1280_nl;
  wire[15:0] Accum2_acc_1274_nl;
  wire[16:0] nl_Accum2_acc_1274_nl;
  wire[19:0] Product1_10_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1273_nl;
  wire[16:0] nl_Accum2_acc_1273_nl;
  wire[19:0] Product1_12_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1279_nl;
  wire[16:0] nl_Accum2_acc_1279_nl;
  wire[9:0] Accum2_acc_1880_nl;
  wire[10:0] nl_Accum2_acc_1880_nl;
  wire[19:0] Product1_1_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1297_nl;
  wire[17:0] nl_Accum2_acc_1297_nl;
  wire[15:0] Accum2_acc_1291_nl;
  wire[16:0] nl_Accum2_acc_1291_nl;
  wire[19:0] Product1_2_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1290_nl;
  wire[16:0] nl_Accum2_acc_1290_nl;
  wire[19:0] Product1_4_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1289_nl;
  wire[16:0] nl_Accum2_acc_1289_nl;
  wire[19:0] Product1_6_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1288_nl;
  wire[16:0] nl_Accum2_acc_1288_nl;
  wire[19:0] Product1_8_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1296_nl;
  wire[16:0] nl_Accum2_acc_1296_nl;
  wire[15:0] Accum2_acc_1293_nl;
  wire[16:0] nl_Accum2_acc_1293_nl;
  wire[15:0] Accum2_acc_1287_nl;
  wire[16:0] nl_Accum2_acc_1287_nl;
  wire[19:0] Product1_10_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1286_nl;
  wire[16:0] nl_Accum2_acc_1286_nl;
  wire[19:0] Product1_12_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1292_nl;
  wire[16:0] nl_Accum2_acc_1292_nl;
  wire[9:0] Accum2_acc_1881_nl;
  wire[10:0] nl_Accum2_acc_1881_nl;
  wire[19:0] Product1_1_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1310_nl;
  wire[17:0] nl_Accum2_acc_1310_nl;
  wire[15:0] Accum2_acc_1304_nl;
  wire[16:0] nl_Accum2_acc_1304_nl;
  wire[19:0] Product1_2_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1303_nl;
  wire[16:0] nl_Accum2_acc_1303_nl;
  wire[19:0] Product1_4_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1302_nl;
  wire[16:0] nl_Accum2_acc_1302_nl;
  wire[19:0] Product1_6_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1301_nl;
  wire[16:0] nl_Accum2_acc_1301_nl;
  wire[19:0] Product1_8_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1309_nl;
  wire[16:0] nl_Accum2_acc_1309_nl;
  wire[15:0] Accum2_acc_1306_nl;
  wire[16:0] nl_Accum2_acc_1306_nl;
  wire[15:0] Accum2_acc_1300_nl;
  wire[16:0] nl_Accum2_acc_1300_nl;
  wire[19:0] Product1_10_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1299_nl;
  wire[16:0] nl_Accum2_acc_1299_nl;
  wire[19:0] Product1_12_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1305_nl;
  wire[16:0] nl_Accum2_acc_1305_nl;
  wire[9:0] Accum2_acc_1882_nl;
  wire[10:0] nl_Accum2_acc_1882_nl;
  wire[19:0] Product1_1_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1323_nl;
  wire[17:0] nl_Accum2_acc_1323_nl;
  wire[15:0] Accum2_acc_1317_nl;
  wire[16:0] nl_Accum2_acc_1317_nl;
  wire[19:0] Product1_2_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1316_nl;
  wire[16:0] nl_Accum2_acc_1316_nl;
  wire[19:0] Product1_4_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1315_nl;
  wire[16:0] nl_Accum2_acc_1315_nl;
  wire[19:0] Product1_6_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1314_nl;
  wire[16:0] nl_Accum2_acc_1314_nl;
  wire[19:0] Product1_8_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1322_nl;
  wire[16:0] nl_Accum2_acc_1322_nl;
  wire[15:0] Accum2_acc_1319_nl;
  wire[16:0] nl_Accum2_acc_1319_nl;
  wire[15:0] Accum2_acc_1313_nl;
  wire[16:0] nl_Accum2_acc_1313_nl;
  wire[19:0] Product1_10_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1312_nl;
  wire[16:0] nl_Accum2_acc_1312_nl;
  wire[19:0] Product1_12_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1318_nl;
  wire[16:0] nl_Accum2_acc_1318_nl;
  wire[9:0] Accum2_acc_1883_nl;
  wire[10:0] nl_Accum2_acc_1883_nl;
  wire[19:0] Product1_1_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1336_nl;
  wire[17:0] nl_Accum2_acc_1336_nl;
  wire[15:0] Accum2_acc_1330_nl;
  wire[16:0] nl_Accum2_acc_1330_nl;
  wire[19:0] Product1_2_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1329_nl;
  wire[16:0] nl_Accum2_acc_1329_nl;
  wire[19:0] Product1_4_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1328_nl;
  wire[16:0] nl_Accum2_acc_1328_nl;
  wire[19:0] Product1_6_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1327_nl;
  wire[16:0] nl_Accum2_acc_1327_nl;
  wire[19:0] Product1_8_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1335_nl;
  wire[16:0] nl_Accum2_acc_1335_nl;
  wire[15:0] Accum2_acc_1332_nl;
  wire[16:0] nl_Accum2_acc_1332_nl;
  wire[15:0] Accum2_acc_1326_nl;
  wire[16:0] nl_Accum2_acc_1326_nl;
  wire[19:0] Product1_10_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1325_nl;
  wire[16:0] nl_Accum2_acc_1325_nl;
  wire[19:0] Product1_12_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1331_nl;
  wire[16:0] nl_Accum2_acc_1331_nl;
  wire[9:0] Accum2_acc_1884_nl;
  wire[10:0] nl_Accum2_acc_1884_nl;
  wire[19:0] Product1_1_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1349_nl;
  wire[17:0] nl_Accum2_acc_1349_nl;
  wire[15:0] Accum2_acc_1343_nl;
  wire[16:0] nl_Accum2_acc_1343_nl;
  wire[19:0] Product1_2_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1342_nl;
  wire[16:0] nl_Accum2_acc_1342_nl;
  wire[19:0] Product1_4_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1341_nl;
  wire[16:0] nl_Accum2_acc_1341_nl;
  wire[19:0] Product1_6_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1340_nl;
  wire[16:0] nl_Accum2_acc_1340_nl;
  wire[19:0] Product1_8_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1348_nl;
  wire[16:0] nl_Accum2_acc_1348_nl;
  wire[15:0] Accum2_acc_1345_nl;
  wire[16:0] nl_Accum2_acc_1345_nl;
  wire[15:0] Accum2_acc_1339_nl;
  wire[16:0] nl_Accum2_acc_1339_nl;
  wire[19:0] Product1_10_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1338_nl;
  wire[16:0] nl_Accum2_acc_1338_nl;
  wire[19:0] Product1_12_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1344_nl;
  wire[16:0] nl_Accum2_acc_1344_nl;
  wire[9:0] Accum2_acc_1885_nl;
  wire[10:0] nl_Accum2_acc_1885_nl;
  wire[19:0] Product1_1_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1362_nl;
  wire[17:0] nl_Accum2_acc_1362_nl;
  wire[15:0] Accum2_acc_1356_nl;
  wire[16:0] nl_Accum2_acc_1356_nl;
  wire[19:0] Product1_2_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1355_nl;
  wire[16:0] nl_Accum2_acc_1355_nl;
  wire[19:0] Product1_4_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1354_nl;
  wire[16:0] nl_Accum2_acc_1354_nl;
  wire[19:0] Product1_6_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1353_nl;
  wire[16:0] nl_Accum2_acc_1353_nl;
  wire[19:0] Product1_8_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1361_nl;
  wire[16:0] nl_Accum2_acc_1361_nl;
  wire[15:0] Accum2_acc_1358_nl;
  wire[16:0] nl_Accum2_acc_1358_nl;
  wire[15:0] Accum2_acc_1352_nl;
  wire[16:0] nl_Accum2_acc_1352_nl;
  wire[19:0] Product1_10_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1351_nl;
  wire[16:0] nl_Accum2_acc_1351_nl;
  wire[19:0] Product1_12_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1357_nl;
  wire[16:0] nl_Accum2_acc_1357_nl;
  wire[9:0] Accum2_acc_1886_nl;
  wire[10:0] nl_Accum2_acc_1886_nl;
  wire[19:0] Product1_1_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1375_nl;
  wire[17:0] nl_Accum2_acc_1375_nl;
  wire[15:0] Accum2_acc_1369_nl;
  wire[16:0] nl_Accum2_acc_1369_nl;
  wire[19:0] Product1_2_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1368_nl;
  wire[16:0] nl_Accum2_acc_1368_nl;
  wire[19:0] Product1_4_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1367_nl;
  wire[16:0] nl_Accum2_acc_1367_nl;
  wire[19:0] Product1_6_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1366_nl;
  wire[16:0] nl_Accum2_acc_1366_nl;
  wire[19:0] Product1_8_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1374_nl;
  wire[16:0] nl_Accum2_acc_1374_nl;
  wire[15:0] Accum2_acc_1371_nl;
  wire[16:0] nl_Accum2_acc_1371_nl;
  wire[15:0] Accum2_acc_1365_nl;
  wire[16:0] nl_Accum2_acc_1365_nl;
  wire[19:0] Product1_10_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1364_nl;
  wire[16:0] nl_Accum2_acc_1364_nl;
  wire[19:0] Product1_12_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1370_nl;
  wire[16:0] nl_Accum2_acc_1370_nl;
  wire[9:0] Accum2_acc_1887_nl;
  wire[10:0] nl_Accum2_acc_1887_nl;
  wire[19:0] Product1_1_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1388_nl;
  wire[17:0] nl_Accum2_acc_1388_nl;
  wire[15:0] Accum2_acc_1382_nl;
  wire[16:0] nl_Accum2_acc_1382_nl;
  wire[19:0] Product1_2_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1381_nl;
  wire[16:0] nl_Accum2_acc_1381_nl;
  wire[19:0] Product1_4_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1380_nl;
  wire[16:0] nl_Accum2_acc_1380_nl;
  wire[19:0] Product1_6_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1379_nl;
  wire[16:0] nl_Accum2_acc_1379_nl;
  wire[19:0] Product1_8_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1387_nl;
  wire[16:0] nl_Accum2_acc_1387_nl;
  wire[15:0] Accum2_acc_1384_nl;
  wire[16:0] nl_Accum2_acc_1384_nl;
  wire[15:0] Accum2_acc_1378_nl;
  wire[16:0] nl_Accum2_acc_1378_nl;
  wire[19:0] Product1_10_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1377_nl;
  wire[16:0] nl_Accum2_acc_1377_nl;
  wire[19:0] Product1_12_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1383_nl;
  wire[16:0] nl_Accum2_acc_1383_nl;
  wire[9:0] Accum2_acc_1888_nl;
  wire[10:0] nl_Accum2_acc_1888_nl;
  wire[19:0] Product1_1_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1401_nl;
  wire[17:0] nl_Accum2_acc_1401_nl;
  wire[15:0] Accum2_acc_1395_nl;
  wire[16:0] nl_Accum2_acc_1395_nl;
  wire[19:0] Product1_2_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1394_nl;
  wire[16:0] nl_Accum2_acc_1394_nl;
  wire[19:0] Product1_4_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1393_nl;
  wire[16:0] nl_Accum2_acc_1393_nl;
  wire[19:0] Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1392_nl;
  wire[16:0] nl_Accum2_acc_1392_nl;
  wire[19:0] Product1_8_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1400_nl;
  wire[16:0] nl_Accum2_acc_1400_nl;
  wire[15:0] Accum2_acc_1397_nl;
  wire[16:0] nl_Accum2_acc_1397_nl;
  wire[15:0] Accum2_acc_1391_nl;
  wire[16:0] nl_Accum2_acc_1391_nl;
  wire[19:0] Product1_10_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1390_nl;
  wire[16:0] nl_Accum2_acc_1390_nl;
  wire[19:0] Product1_12_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1396_nl;
  wire[16:0] nl_Accum2_acc_1396_nl;
  wire[9:0] Accum2_acc_1889_nl;
  wire[10:0] nl_Accum2_acc_1889_nl;
  wire[19:0] Product1_1_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1414_nl;
  wire[17:0] nl_Accum2_acc_1414_nl;
  wire[15:0] Accum2_acc_1408_nl;
  wire[16:0] nl_Accum2_acc_1408_nl;
  wire[19:0] Product1_2_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1407_nl;
  wire[16:0] nl_Accum2_acc_1407_nl;
  wire[19:0] Product1_4_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1406_nl;
  wire[16:0] nl_Accum2_acc_1406_nl;
  wire[19:0] Product1_6_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1405_nl;
  wire[16:0] nl_Accum2_acc_1405_nl;
  wire[19:0] Product1_8_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1413_nl;
  wire[16:0] nl_Accum2_acc_1413_nl;
  wire[15:0] Accum2_acc_1410_nl;
  wire[16:0] nl_Accum2_acc_1410_nl;
  wire[15:0] Accum2_acc_1404_nl;
  wire[16:0] nl_Accum2_acc_1404_nl;
  wire[19:0] Product1_10_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1403_nl;
  wire[16:0] nl_Accum2_acc_1403_nl;
  wire[19:0] Product1_12_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1409_nl;
  wire[16:0] nl_Accum2_acc_1409_nl;
  wire[9:0] Accum2_acc_1890_nl;
  wire[10:0] nl_Accum2_acc_1890_nl;
  wire[19:0] Product1_1_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1427_nl;
  wire[17:0] nl_Accum2_acc_1427_nl;
  wire[15:0] Accum2_acc_1421_nl;
  wire[16:0] nl_Accum2_acc_1421_nl;
  wire[19:0] Product1_2_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1420_nl;
  wire[16:0] nl_Accum2_acc_1420_nl;
  wire[19:0] Product1_4_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1419_nl;
  wire[16:0] nl_Accum2_acc_1419_nl;
  wire[19:0] Product1_6_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1418_nl;
  wire[16:0] nl_Accum2_acc_1418_nl;
  wire[19:0] Product1_8_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1426_nl;
  wire[16:0] nl_Accum2_acc_1426_nl;
  wire[15:0] Accum2_acc_1423_nl;
  wire[16:0] nl_Accum2_acc_1423_nl;
  wire[15:0] Accum2_acc_1417_nl;
  wire[16:0] nl_Accum2_acc_1417_nl;
  wire[19:0] Product1_10_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1416_nl;
  wire[16:0] nl_Accum2_acc_1416_nl;
  wire[19:0] Product1_12_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1422_nl;
  wire[16:0] nl_Accum2_acc_1422_nl;
  wire[9:0] Accum2_acc_1891_nl;
  wire[10:0] nl_Accum2_acc_1891_nl;
  wire[19:0] Product1_1_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1440_nl;
  wire[17:0] nl_Accum2_acc_1440_nl;
  wire[15:0] Accum2_acc_1434_nl;
  wire[16:0] nl_Accum2_acc_1434_nl;
  wire[19:0] Product1_2_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1433_nl;
  wire[16:0] nl_Accum2_acc_1433_nl;
  wire[19:0] Product1_4_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1432_nl;
  wire[16:0] nl_Accum2_acc_1432_nl;
  wire[19:0] Product1_6_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1431_nl;
  wire[16:0] nl_Accum2_acc_1431_nl;
  wire[19:0] Product1_8_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1439_nl;
  wire[16:0] nl_Accum2_acc_1439_nl;
  wire[15:0] Accum2_acc_1436_nl;
  wire[16:0] nl_Accum2_acc_1436_nl;
  wire[15:0] Accum2_acc_1430_nl;
  wire[16:0] nl_Accum2_acc_1430_nl;
  wire[19:0] Product1_10_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1429_nl;
  wire[16:0] nl_Accum2_acc_1429_nl;
  wire[19:0] Product1_12_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1435_nl;
  wire[16:0] nl_Accum2_acc_1435_nl;
  wire[9:0] Accum2_acc_1892_nl;
  wire[10:0] nl_Accum2_acc_1892_nl;
  wire[19:0] Product1_1_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1453_nl;
  wire[17:0] nl_Accum2_acc_1453_nl;
  wire[15:0] Accum2_acc_1447_nl;
  wire[16:0] nl_Accum2_acc_1447_nl;
  wire[19:0] Product1_2_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1446_nl;
  wire[16:0] nl_Accum2_acc_1446_nl;
  wire[19:0] Product1_4_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1445_nl;
  wire[16:0] nl_Accum2_acc_1445_nl;
  wire[19:0] Product1_6_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1444_nl;
  wire[16:0] nl_Accum2_acc_1444_nl;
  wire[19:0] Product1_8_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1452_nl;
  wire[16:0] nl_Accum2_acc_1452_nl;
  wire[15:0] Accum2_acc_1449_nl;
  wire[16:0] nl_Accum2_acc_1449_nl;
  wire[15:0] Accum2_acc_1443_nl;
  wire[16:0] nl_Accum2_acc_1443_nl;
  wire[19:0] Product1_10_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1442_nl;
  wire[16:0] nl_Accum2_acc_1442_nl;
  wire[19:0] Product1_12_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1448_nl;
  wire[16:0] nl_Accum2_acc_1448_nl;
  wire[9:0] Accum2_acc_1893_nl;
  wire[10:0] nl_Accum2_acc_1893_nl;
  wire[19:0] Product1_1_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1466_nl;
  wire[17:0] nl_Accum2_acc_1466_nl;
  wire[15:0] Accum2_acc_1460_nl;
  wire[16:0] nl_Accum2_acc_1460_nl;
  wire[19:0] Product1_2_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1459_nl;
  wire[16:0] nl_Accum2_acc_1459_nl;
  wire[19:0] Product1_4_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1458_nl;
  wire[16:0] nl_Accum2_acc_1458_nl;
  wire[19:0] Product1_6_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1457_nl;
  wire[16:0] nl_Accum2_acc_1457_nl;
  wire[19:0] Product1_8_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1465_nl;
  wire[16:0] nl_Accum2_acc_1465_nl;
  wire[15:0] Accum2_acc_1462_nl;
  wire[16:0] nl_Accum2_acc_1462_nl;
  wire[15:0] Accum2_acc_1456_nl;
  wire[16:0] nl_Accum2_acc_1456_nl;
  wire[19:0] Product1_10_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1455_nl;
  wire[16:0] nl_Accum2_acc_1455_nl;
  wire[19:0] Product1_12_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1461_nl;
  wire[16:0] nl_Accum2_acc_1461_nl;
  wire[9:0] Accum2_acc_1894_nl;
  wire[10:0] nl_Accum2_acc_1894_nl;
  wire[19:0] Product1_1_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1479_nl;
  wire[17:0] nl_Accum2_acc_1479_nl;
  wire[15:0] Accum2_acc_1473_nl;
  wire[16:0] nl_Accum2_acc_1473_nl;
  wire[19:0] Product1_2_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1472_nl;
  wire[16:0] nl_Accum2_acc_1472_nl;
  wire[19:0] Product1_4_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1471_nl;
  wire[16:0] nl_Accum2_acc_1471_nl;
  wire[19:0] Product1_6_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1470_nl;
  wire[16:0] nl_Accum2_acc_1470_nl;
  wire[19:0] Product1_8_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1478_nl;
  wire[16:0] nl_Accum2_acc_1478_nl;
  wire[15:0] Accum2_acc_1475_nl;
  wire[16:0] nl_Accum2_acc_1475_nl;
  wire[15:0] Accum2_acc_1469_nl;
  wire[16:0] nl_Accum2_acc_1469_nl;
  wire[19:0] Product1_10_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1468_nl;
  wire[16:0] nl_Accum2_acc_1468_nl;
  wire[19:0] Product1_12_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1474_nl;
  wire[16:0] nl_Accum2_acc_1474_nl;
  wire[9:0] Accum2_acc_1895_nl;
  wire[10:0] nl_Accum2_acc_1895_nl;
  wire[19:0] Product1_1_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1492_nl;
  wire[17:0] nl_Accum2_acc_1492_nl;
  wire[15:0] Accum2_acc_1486_nl;
  wire[16:0] nl_Accum2_acc_1486_nl;
  wire[19:0] Product1_2_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1485_nl;
  wire[16:0] nl_Accum2_acc_1485_nl;
  wire[19:0] Product1_4_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1484_nl;
  wire[16:0] nl_Accum2_acc_1484_nl;
  wire[19:0] Product1_6_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1483_nl;
  wire[16:0] nl_Accum2_acc_1483_nl;
  wire[19:0] Product1_8_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1491_nl;
  wire[16:0] nl_Accum2_acc_1491_nl;
  wire[15:0] Accum2_acc_1488_nl;
  wire[16:0] nl_Accum2_acc_1488_nl;
  wire[15:0] Accum2_acc_1482_nl;
  wire[16:0] nl_Accum2_acc_1482_nl;
  wire[19:0] Product1_10_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1481_nl;
  wire[16:0] nl_Accum2_acc_1481_nl;
  wire[19:0] Product1_12_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1487_nl;
  wire[16:0] nl_Accum2_acc_1487_nl;
  wire[9:0] Accum2_acc_1896_nl;
  wire[10:0] nl_Accum2_acc_1896_nl;
  wire[19:0] Product1_1_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1505_nl;
  wire[17:0] nl_Accum2_acc_1505_nl;
  wire[15:0] Accum2_acc_1499_nl;
  wire[16:0] nl_Accum2_acc_1499_nl;
  wire[19:0] Product1_2_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1498_nl;
  wire[16:0] nl_Accum2_acc_1498_nl;
  wire[19:0] Product1_4_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1497_nl;
  wire[16:0] nl_Accum2_acc_1497_nl;
  wire[19:0] Product1_6_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1496_nl;
  wire[16:0] nl_Accum2_acc_1496_nl;
  wire[19:0] Product1_8_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1504_nl;
  wire[16:0] nl_Accum2_acc_1504_nl;
  wire[15:0] Accum2_acc_1501_nl;
  wire[16:0] nl_Accum2_acc_1501_nl;
  wire[15:0] Accum2_acc_1495_nl;
  wire[16:0] nl_Accum2_acc_1495_nl;
  wire[19:0] Product1_10_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1494_nl;
  wire[16:0] nl_Accum2_acc_1494_nl;
  wire[19:0] Product1_12_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1500_nl;
  wire[16:0] nl_Accum2_acc_1500_nl;
  wire[9:0] Accum2_acc_1897_nl;
  wire[10:0] nl_Accum2_acc_1897_nl;
  wire[19:0] Product1_1_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1518_nl;
  wire[17:0] nl_Accum2_acc_1518_nl;
  wire[15:0] Accum2_acc_1512_nl;
  wire[16:0] nl_Accum2_acc_1512_nl;
  wire[19:0] Product1_2_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1511_nl;
  wire[16:0] nl_Accum2_acc_1511_nl;
  wire[19:0] Product1_4_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1510_nl;
  wire[16:0] nl_Accum2_acc_1510_nl;
  wire[19:0] Product1_6_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1509_nl;
  wire[16:0] nl_Accum2_acc_1509_nl;
  wire[19:0] Product1_8_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1517_nl;
  wire[16:0] nl_Accum2_acc_1517_nl;
  wire[15:0] Accum2_acc_1514_nl;
  wire[16:0] nl_Accum2_acc_1514_nl;
  wire[15:0] Accum2_acc_1508_nl;
  wire[16:0] nl_Accum2_acc_1508_nl;
  wire[19:0] Product1_10_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1507_nl;
  wire[16:0] nl_Accum2_acc_1507_nl;
  wire[19:0] Product1_12_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1513_nl;
  wire[16:0] nl_Accum2_acc_1513_nl;
  wire[9:0] Accum2_acc_1898_nl;
  wire[10:0] nl_Accum2_acc_1898_nl;
  wire[19:0] Product1_1_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1531_nl;
  wire[17:0] nl_Accum2_acc_1531_nl;
  wire[15:0] Accum2_acc_1525_nl;
  wire[16:0] nl_Accum2_acc_1525_nl;
  wire[19:0] Product1_2_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1524_nl;
  wire[16:0] nl_Accum2_acc_1524_nl;
  wire[19:0] Product1_4_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1523_nl;
  wire[16:0] nl_Accum2_acc_1523_nl;
  wire[19:0] Product1_6_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1522_nl;
  wire[16:0] nl_Accum2_acc_1522_nl;
  wire[19:0] Product1_8_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1530_nl;
  wire[16:0] nl_Accum2_acc_1530_nl;
  wire[15:0] Accum2_acc_1527_nl;
  wire[16:0] nl_Accum2_acc_1527_nl;
  wire[15:0] Accum2_acc_1521_nl;
  wire[16:0] nl_Accum2_acc_1521_nl;
  wire[19:0] Product1_10_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1520_nl;
  wire[16:0] nl_Accum2_acc_1520_nl;
  wire[19:0] Product1_12_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1526_nl;
  wire[16:0] nl_Accum2_acc_1526_nl;
  wire[9:0] Accum2_acc_1899_nl;
  wire[10:0] nl_Accum2_acc_1899_nl;
  wire[19:0] Product1_1_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1544_nl;
  wire[17:0] nl_Accum2_acc_1544_nl;
  wire[15:0] Accum2_acc_1538_nl;
  wire[16:0] nl_Accum2_acc_1538_nl;
  wire[19:0] Product1_2_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1537_nl;
  wire[16:0] nl_Accum2_acc_1537_nl;
  wire[19:0] Product1_4_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1536_nl;
  wire[16:0] nl_Accum2_acc_1536_nl;
  wire[19:0] Product1_6_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1535_nl;
  wire[16:0] nl_Accum2_acc_1535_nl;
  wire[19:0] Product1_8_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1543_nl;
  wire[16:0] nl_Accum2_acc_1543_nl;
  wire[15:0] Accum2_acc_1540_nl;
  wire[16:0] nl_Accum2_acc_1540_nl;
  wire[15:0] Accum2_acc_1534_nl;
  wire[16:0] nl_Accum2_acc_1534_nl;
  wire[19:0] Product1_10_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1533_nl;
  wire[16:0] nl_Accum2_acc_1533_nl;
  wire[19:0] Product1_12_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1539_nl;
  wire[16:0] nl_Accum2_acc_1539_nl;
  wire[9:0] Accum2_acc_1900_nl;
  wire[10:0] nl_Accum2_acc_1900_nl;
  wire[19:0] Product1_1_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1557_nl;
  wire[17:0] nl_Accum2_acc_1557_nl;
  wire[15:0] Accum2_acc_1551_nl;
  wire[16:0] nl_Accum2_acc_1551_nl;
  wire[19:0] Product1_2_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1550_nl;
  wire[16:0] nl_Accum2_acc_1550_nl;
  wire[19:0] Product1_4_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1549_nl;
  wire[16:0] nl_Accum2_acc_1549_nl;
  wire[19:0] Product1_6_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1548_nl;
  wire[16:0] nl_Accum2_acc_1548_nl;
  wire[19:0] Product1_8_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1556_nl;
  wire[16:0] nl_Accum2_acc_1556_nl;
  wire[15:0] Accum2_acc_1553_nl;
  wire[16:0] nl_Accum2_acc_1553_nl;
  wire[15:0] Accum2_acc_1547_nl;
  wire[16:0] nl_Accum2_acc_1547_nl;
  wire[19:0] Product1_10_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1546_nl;
  wire[16:0] nl_Accum2_acc_1546_nl;
  wire[19:0] Product1_12_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1552_nl;
  wire[16:0] nl_Accum2_acc_1552_nl;
  wire[9:0] Accum2_acc_1901_nl;
  wire[10:0] nl_Accum2_acc_1901_nl;
  wire[19:0] Product1_1_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1570_nl;
  wire[17:0] nl_Accum2_acc_1570_nl;
  wire[15:0] Accum2_acc_1564_nl;
  wire[16:0] nl_Accum2_acc_1564_nl;
  wire[19:0] Product1_2_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1563_nl;
  wire[16:0] nl_Accum2_acc_1563_nl;
  wire[19:0] Product1_4_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1562_nl;
  wire[16:0] nl_Accum2_acc_1562_nl;
  wire[19:0] Product1_6_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1561_nl;
  wire[16:0] nl_Accum2_acc_1561_nl;
  wire[19:0] Product1_8_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1569_nl;
  wire[16:0] nl_Accum2_acc_1569_nl;
  wire[15:0] Accum2_acc_1566_nl;
  wire[16:0] nl_Accum2_acc_1566_nl;
  wire[15:0] Accum2_acc_1560_nl;
  wire[16:0] nl_Accum2_acc_1560_nl;
  wire[19:0] Product1_10_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1559_nl;
  wire[16:0] nl_Accum2_acc_1559_nl;
  wire[19:0] Product1_12_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1565_nl;
  wire[16:0] nl_Accum2_acc_1565_nl;
  wire[9:0] Accum2_acc_1902_nl;
  wire[10:0] nl_Accum2_acc_1902_nl;
  wire[19:0] Product1_1_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1583_nl;
  wire[17:0] nl_Accum2_acc_1583_nl;
  wire[15:0] Accum2_acc_1577_nl;
  wire[16:0] nl_Accum2_acc_1577_nl;
  wire[19:0] Product1_2_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1576_nl;
  wire[16:0] nl_Accum2_acc_1576_nl;
  wire[19:0] Product1_4_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1575_nl;
  wire[16:0] nl_Accum2_acc_1575_nl;
  wire[19:0] Product1_6_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1574_nl;
  wire[16:0] nl_Accum2_acc_1574_nl;
  wire[19:0] Product1_8_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1582_nl;
  wire[16:0] nl_Accum2_acc_1582_nl;
  wire[15:0] Accum2_acc_1579_nl;
  wire[16:0] nl_Accum2_acc_1579_nl;
  wire[15:0] Accum2_acc_1573_nl;
  wire[16:0] nl_Accum2_acc_1573_nl;
  wire[19:0] Product1_10_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1572_nl;
  wire[16:0] nl_Accum2_acc_1572_nl;
  wire[19:0] Product1_12_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1578_nl;
  wire[16:0] nl_Accum2_acc_1578_nl;
  wire[9:0] Accum2_acc_1903_nl;
  wire[10:0] nl_Accum2_acc_1903_nl;
  wire[19:0] Product1_1_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1596_nl;
  wire[17:0] nl_Accum2_acc_1596_nl;
  wire[15:0] Accum2_acc_1590_nl;
  wire[16:0] nl_Accum2_acc_1590_nl;
  wire[19:0] Product1_2_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1589_nl;
  wire[16:0] nl_Accum2_acc_1589_nl;
  wire[19:0] Product1_4_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1588_nl;
  wire[16:0] nl_Accum2_acc_1588_nl;
  wire[19:0] Product1_6_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1587_nl;
  wire[16:0] nl_Accum2_acc_1587_nl;
  wire[19:0] Product1_8_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1595_nl;
  wire[16:0] nl_Accum2_acc_1595_nl;
  wire[15:0] Accum2_acc_1592_nl;
  wire[16:0] nl_Accum2_acc_1592_nl;
  wire[15:0] Accum2_acc_1586_nl;
  wire[16:0] nl_Accum2_acc_1586_nl;
  wire[19:0] Product1_10_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1585_nl;
  wire[16:0] nl_Accum2_acc_1585_nl;
  wire[19:0] Product1_12_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1591_nl;
  wire[16:0] nl_Accum2_acc_1591_nl;
  wire[9:0] Accum2_acc_1904_nl;
  wire[10:0] nl_Accum2_acc_1904_nl;
  wire[19:0] Product1_1_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1609_nl;
  wire[17:0] nl_Accum2_acc_1609_nl;
  wire[15:0] Accum2_acc_1603_nl;
  wire[16:0] nl_Accum2_acc_1603_nl;
  wire[19:0] Product1_2_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1602_nl;
  wire[16:0] nl_Accum2_acc_1602_nl;
  wire[19:0] Product1_4_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1601_nl;
  wire[16:0] nl_Accum2_acc_1601_nl;
  wire[19:0] Product1_6_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1600_nl;
  wire[16:0] nl_Accum2_acc_1600_nl;
  wire[19:0] Product1_8_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1608_nl;
  wire[16:0] nl_Accum2_acc_1608_nl;
  wire[15:0] Accum2_acc_1605_nl;
  wire[16:0] nl_Accum2_acc_1605_nl;
  wire[15:0] Accum2_acc_1599_nl;
  wire[16:0] nl_Accum2_acc_1599_nl;
  wire[19:0] Product1_10_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1598_nl;
  wire[16:0] nl_Accum2_acc_1598_nl;
  wire[19:0] Product1_12_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1604_nl;
  wire[16:0] nl_Accum2_acc_1604_nl;
  wire[9:0] Accum2_acc_1905_nl;
  wire[10:0] nl_Accum2_acc_1905_nl;
  wire[19:0] Product1_1_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1622_nl;
  wire[17:0] nl_Accum2_acc_1622_nl;
  wire[15:0] Accum2_acc_1616_nl;
  wire[16:0] nl_Accum2_acc_1616_nl;
  wire[19:0] Product1_2_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1615_nl;
  wire[16:0] nl_Accum2_acc_1615_nl;
  wire[19:0] Product1_4_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1614_nl;
  wire[16:0] nl_Accum2_acc_1614_nl;
  wire[19:0] Product1_6_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1613_nl;
  wire[16:0] nl_Accum2_acc_1613_nl;
  wire[19:0] Product1_8_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1621_nl;
  wire[16:0] nl_Accum2_acc_1621_nl;
  wire[15:0] Accum2_acc_1618_nl;
  wire[16:0] nl_Accum2_acc_1618_nl;
  wire[15:0] Accum2_acc_1612_nl;
  wire[16:0] nl_Accum2_acc_1612_nl;
  wire[19:0] Product1_10_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1611_nl;
  wire[16:0] nl_Accum2_acc_1611_nl;
  wire[19:0] Product1_12_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1617_nl;
  wire[16:0] nl_Accum2_acc_1617_nl;
  wire[9:0] Accum2_acc_1906_nl;
  wire[10:0] nl_Accum2_acc_1906_nl;
  wire[19:0] Product1_1_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1635_nl;
  wire[17:0] nl_Accum2_acc_1635_nl;
  wire[15:0] Accum2_acc_1629_nl;
  wire[16:0] nl_Accum2_acc_1629_nl;
  wire[19:0] Product1_2_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1628_nl;
  wire[16:0] nl_Accum2_acc_1628_nl;
  wire[19:0] Product1_4_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1627_nl;
  wire[16:0] nl_Accum2_acc_1627_nl;
  wire[19:0] Product1_6_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1626_nl;
  wire[16:0] nl_Accum2_acc_1626_nl;
  wire[19:0] Product1_8_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1634_nl;
  wire[16:0] nl_Accum2_acc_1634_nl;
  wire[15:0] Accum2_acc_1631_nl;
  wire[16:0] nl_Accum2_acc_1631_nl;
  wire[15:0] Accum2_acc_1625_nl;
  wire[16:0] nl_Accum2_acc_1625_nl;
  wire[19:0] Product1_10_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1624_nl;
  wire[16:0] nl_Accum2_acc_1624_nl;
  wire[19:0] Product1_12_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1630_nl;
  wire[16:0] nl_Accum2_acc_1630_nl;
  wire[9:0] Accum2_acc_1907_nl;
  wire[10:0] nl_Accum2_acc_1907_nl;
  wire[19:0] Product1_1_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1648_nl;
  wire[17:0] nl_Accum2_acc_1648_nl;
  wire[15:0] Accum2_acc_1642_nl;
  wire[16:0] nl_Accum2_acc_1642_nl;
  wire[19:0] Product1_2_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1641_nl;
  wire[16:0] nl_Accum2_acc_1641_nl;
  wire[19:0] Product1_4_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1640_nl;
  wire[16:0] nl_Accum2_acc_1640_nl;
  wire[19:0] Product1_6_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1639_nl;
  wire[16:0] nl_Accum2_acc_1639_nl;
  wire[19:0] Product1_8_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1647_nl;
  wire[16:0] nl_Accum2_acc_1647_nl;
  wire[15:0] Accum2_acc_1644_nl;
  wire[16:0] nl_Accum2_acc_1644_nl;
  wire[15:0] Accum2_acc_1638_nl;
  wire[16:0] nl_Accum2_acc_1638_nl;
  wire[19:0] Product1_10_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1637_nl;
  wire[16:0] nl_Accum2_acc_1637_nl;
  wire[19:0] Product1_12_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1643_nl;
  wire[16:0] nl_Accum2_acc_1643_nl;
  wire[9:0] Accum2_acc_1908_nl;
  wire[10:0] nl_Accum2_acc_1908_nl;
  wire[19:0] Product1_1_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1661_nl;
  wire[17:0] nl_Accum2_acc_1661_nl;
  wire[15:0] Accum2_acc_1655_nl;
  wire[16:0] nl_Accum2_acc_1655_nl;
  wire[19:0] Product1_2_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1654_nl;
  wire[16:0] nl_Accum2_acc_1654_nl;
  wire[19:0] Product1_4_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1653_nl;
  wire[16:0] nl_Accum2_acc_1653_nl;
  wire[19:0] Product1_6_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1652_nl;
  wire[16:0] nl_Accum2_acc_1652_nl;
  wire[19:0] Product1_8_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1660_nl;
  wire[16:0] nl_Accum2_acc_1660_nl;
  wire[15:0] Accum2_acc_1657_nl;
  wire[16:0] nl_Accum2_acc_1657_nl;
  wire[15:0] Accum2_acc_1651_nl;
  wire[16:0] nl_Accum2_acc_1651_nl;
  wire[19:0] Product1_10_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1650_nl;
  wire[16:0] nl_Accum2_acc_1650_nl;
  wire[19:0] Product1_12_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1656_nl;
  wire[16:0] nl_Accum2_acc_1656_nl;
  wire[9:0] Accum2_acc_1909_nl;
  wire[10:0] nl_Accum2_acc_1909_nl;
  wire[19:0] Product1_1_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1674_nl;
  wire[17:0] nl_Accum2_acc_1674_nl;
  wire[15:0] Accum2_acc_1668_nl;
  wire[16:0] nl_Accum2_acc_1668_nl;
  wire[19:0] Product1_2_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1667_nl;
  wire[16:0] nl_Accum2_acc_1667_nl;
  wire[19:0] Product1_4_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1666_nl;
  wire[16:0] nl_Accum2_acc_1666_nl;
  wire[19:0] Product1_6_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1665_nl;
  wire[16:0] nl_Accum2_acc_1665_nl;
  wire[19:0] Product1_8_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1673_nl;
  wire[16:0] nl_Accum2_acc_1673_nl;
  wire[15:0] Accum2_acc_1670_nl;
  wire[16:0] nl_Accum2_acc_1670_nl;
  wire[15:0] Accum2_acc_1664_nl;
  wire[16:0] nl_Accum2_acc_1664_nl;
  wire[19:0] Product1_10_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1663_nl;
  wire[16:0] nl_Accum2_acc_1663_nl;
  wire[19:0] Product1_12_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1669_nl;
  wire[16:0] nl_Accum2_acc_1669_nl;
  wire[9:0] Accum2_acc_1910_nl;
  wire[10:0] nl_Accum2_acc_1910_nl;
  wire[19:0] Product1_1_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1687_nl;
  wire[17:0] nl_Accum2_acc_1687_nl;
  wire[15:0] Accum2_acc_1681_nl;
  wire[16:0] nl_Accum2_acc_1681_nl;
  wire[19:0] Product1_2_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1680_nl;
  wire[16:0] nl_Accum2_acc_1680_nl;
  wire[19:0] Product1_4_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1679_nl;
  wire[16:0] nl_Accum2_acc_1679_nl;
  wire[19:0] Product1_6_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1678_nl;
  wire[16:0] nl_Accum2_acc_1678_nl;
  wire[19:0] Product1_8_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1686_nl;
  wire[16:0] nl_Accum2_acc_1686_nl;
  wire[15:0] Accum2_acc_1683_nl;
  wire[16:0] nl_Accum2_acc_1683_nl;
  wire[15:0] Accum2_acc_1677_nl;
  wire[16:0] nl_Accum2_acc_1677_nl;
  wire[19:0] Product1_10_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1676_nl;
  wire[16:0] nl_Accum2_acc_1676_nl;
  wire[19:0] Product1_12_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1682_nl;
  wire[16:0] nl_Accum2_acc_1682_nl;
  wire[9:0] Accum2_acc_1911_nl;
  wire[10:0] nl_Accum2_acc_1911_nl;
  wire[19:0] Product1_1_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1700_nl;
  wire[17:0] nl_Accum2_acc_1700_nl;
  wire[15:0] Accum2_acc_1694_nl;
  wire[16:0] nl_Accum2_acc_1694_nl;
  wire[19:0] Product1_2_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1693_nl;
  wire[16:0] nl_Accum2_acc_1693_nl;
  wire[19:0] Product1_4_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1692_nl;
  wire[16:0] nl_Accum2_acc_1692_nl;
  wire[19:0] Product1_6_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1691_nl;
  wire[16:0] nl_Accum2_acc_1691_nl;
  wire[19:0] Product1_8_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1699_nl;
  wire[16:0] nl_Accum2_acc_1699_nl;
  wire[15:0] Accum2_acc_1696_nl;
  wire[16:0] nl_Accum2_acc_1696_nl;
  wire[15:0] Accum2_acc_1690_nl;
  wire[16:0] nl_Accum2_acc_1690_nl;
  wire[19:0] Product1_10_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1689_nl;
  wire[16:0] nl_Accum2_acc_1689_nl;
  wire[19:0] Product1_12_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1695_nl;
  wire[16:0] nl_Accum2_acc_1695_nl;
  wire[9:0] Accum2_acc_1912_nl;
  wire[10:0] nl_Accum2_acc_1912_nl;
  wire[19:0] Product1_1_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1713_nl;
  wire[17:0] nl_Accum2_acc_1713_nl;
  wire[15:0] Accum2_acc_1707_nl;
  wire[16:0] nl_Accum2_acc_1707_nl;
  wire[19:0] Product1_2_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1706_nl;
  wire[16:0] nl_Accum2_acc_1706_nl;
  wire[19:0] Product1_4_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1705_nl;
  wire[16:0] nl_Accum2_acc_1705_nl;
  wire[19:0] Product1_6_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1704_nl;
  wire[16:0] nl_Accum2_acc_1704_nl;
  wire[19:0] Product1_8_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1712_nl;
  wire[16:0] nl_Accum2_acc_1712_nl;
  wire[15:0] Accum2_acc_1709_nl;
  wire[16:0] nl_Accum2_acc_1709_nl;
  wire[15:0] Accum2_acc_1703_nl;
  wire[16:0] nl_Accum2_acc_1703_nl;
  wire[19:0] Product1_10_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1702_nl;
  wire[16:0] nl_Accum2_acc_1702_nl;
  wire[19:0] Product1_12_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1708_nl;
  wire[16:0] nl_Accum2_acc_1708_nl;
  wire[9:0] Accum2_acc_1913_nl;
  wire[10:0] nl_Accum2_acc_1913_nl;
  wire[19:0] Product1_1_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1726_nl;
  wire[17:0] nl_Accum2_acc_1726_nl;
  wire[15:0] Accum2_acc_1720_nl;
  wire[16:0] nl_Accum2_acc_1720_nl;
  wire[19:0] Product1_2_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1719_nl;
  wire[16:0] nl_Accum2_acc_1719_nl;
  wire[19:0] Product1_4_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1718_nl;
  wire[16:0] nl_Accum2_acc_1718_nl;
  wire[19:0] Product1_6_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1717_nl;
  wire[16:0] nl_Accum2_acc_1717_nl;
  wire[19:0] Product1_8_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1725_nl;
  wire[16:0] nl_Accum2_acc_1725_nl;
  wire[15:0] Accum2_acc_1722_nl;
  wire[16:0] nl_Accum2_acc_1722_nl;
  wire[15:0] Accum2_acc_1716_nl;
  wire[16:0] nl_Accum2_acc_1716_nl;
  wire[19:0] Product1_10_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1715_nl;
  wire[16:0] nl_Accum2_acc_1715_nl;
  wire[19:0] Product1_12_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1721_nl;
  wire[16:0] nl_Accum2_acc_1721_nl;
  wire[9:0] Accum2_acc_1914_nl;
  wire[10:0] nl_Accum2_acc_1914_nl;
  wire[19:0] Product1_1_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1739_nl;
  wire[17:0] nl_Accum2_acc_1739_nl;
  wire[15:0] Accum2_acc_1733_nl;
  wire[16:0] nl_Accum2_acc_1733_nl;
  wire[19:0] Product1_2_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1732_nl;
  wire[16:0] nl_Accum2_acc_1732_nl;
  wire[19:0] Product1_4_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1731_nl;
  wire[16:0] nl_Accum2_acc_1731_nl;
  wire[19:0] Product1_6_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1730_nl;
  wire[16:0] nl_Accum2_acc_1730_nl;
  wire[19:0] Product1_8_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1738_nl;
  wire[16:0] nl_Accum2_acc_1738_nl;
  wire[15:0] Accum2_acc_1735_nl;
  wire[16:0] nl_Accum2_acc_1735_nl;
  wire[15:0] Accum2_acc_1729_nl;
  wire[16:0] nl_Accum2_acc_1729_nl;
  wire[19:0] Product1_10_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1728_nl;
  wire[16:0] nl_Accum2_acc_1728_nl;
  wire[19:0] Product1_12_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1734_nl;
  wire[16:0] nl_Accum2_acc_1734_nl;
  wire[9:0] Accum2_acc_1915_nl;
  wire[10:0] nl_Accum2_acc_1915_nl;
  wire[19:0] Product1_1_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1752_nl;
  wire[17:0] nl_Accum2_acc_1752_nl;
  wire[15:0] Accum2_acc_1746_nl;
  wire[16:0] nl_Accum2_acc_1746_nl;
  wire[19:0] Product1_2_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1745_nl;
  wire[16:0] nl_Accum2_acc_1745_nl;
  wire[19:0] Product1_4_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1744_nl;
  wire[16:0] nl_Accum2_acc_1744_nl;
  wire[19:0] Product1_6_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1743_nl;
  wire[16:0] nl_Accum2_acc_1743_nl;
  wire[19:0] Product1_8_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1751_nl;
  wire[16:0] nl_Accum2_acc_1751_nl;
  wire[15:0] Accum2_acc_1748_nl;
  wire[16:0] nl_Accum2_acc_1748_nl;
  wire[15:0] Accum2_acc_1742_nl;
  wire[16:0] nl_Accum2_acc_1742_nl;
  wire[19:0] Product1_10_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1741_nl;
  wire[16:0] nl_Accum2_acc_1741_nl;
  wire[19:0] Product1_12_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1747_nl;
  wire[16:0] nl_Accum2_acc_1747_nl;
  wire[9:0] Accum2_acc_1916_nl;
  wire[10:0] nl_Accum2_acc_1916_nl;
  wire[19:0] Product1_1_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1765_nl;
  wire[17:0] nl_Accum2_acc_1765_nl;
  wire[15:0] Accum2_acc_1759_nl;
  wire[16:0] nl_Accum2_acc_1759_nl;
  wire[19:0] Product1_2_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1758_nl;
  wire[16:0] nl_Accum2_acc_1758_nl;
  wire[19:0] Product1_4_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1757_nl;
  wire[16:0] nl_Accum2_acc_1757_nl;
  wire[19:0] Product1_6_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1756_nl;
  wire[16:0] nl_Accum2_acc_1756_nl;
  wire[19:0] Product1_8_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1764_nl;
  wire[16:0] nl_Accum2_acc_1764_nl;
  wire[15:0] Accum2_acc_1761_nl;
  wire[16:0] nl_Accum2_acc_1761_nl;
  wire[15:0] Accum2_acc_1755_nl;
  wire[16:0] nl_Accum2_acc_1755_nl;
  wire[19:0] Product1_10_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1754_nl;
  wire[16:0] nl_Accum2_acc_1754_nl;
  wire[19:0] Product1_12_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1760_nl;
  wire[16:0] nl_Accum2_acc_1760_nl;
  wire[9:0] Accum2_acc_1917_nl;
  wire[10:0] nl_Accum2_acc_1917_nl;
  wire[19:0] Product1_1_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1778_nl;
  wire[17:0] nl_Accum2_acc_1778_nl;
  wire[15:0] Accum2_acc_1772_nl;
  wire[16:0] nl_Accum2_acc_1772_nl;
  wire[19:0] Product1_2_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1771_nl;
  wire[16:0] nl_Accum2_acc_1771_nl;
  wire[19:0] Product1_4_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1770_nl;
  wire[16:0] nl_Accum2_acc_1770_nl;
  wire[19:0] Product1_6_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1769_nl;
  wire[16:0] nl_Accum2_acc_1769_nl;
  wire[19:0] Product1_8_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1777_nl;
  wire[16:0] nl_Accum2_acc_1777_nl;
  wire[15:0] Accum2_acc_1774_nl;
  wire[16:0] nl_Accum2_acc_1774_nl;
  wire[15:0] Accum2_acc_1768_nl;
  wire[16:0] nl_Accum2_acc_1768_nl;
  wire[19:0] Product1_10_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1767_nl;
  wire[16:0] nl_Accum2_acc_1767_nl;
  wire[19:0] Product1_12_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1773_nl;
  wire[16:0] nl_Accum2_acc_1773_nl;
  wire[9:0] Accum2_acc_1918_nl;
  wire[10:0] nl_Accum2_acc_1918_nl;
  wire[19:0] Product1_1_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1791_nl;
  wire[17:0] nl_Accum2_acc_1791_nl;
  wire[15:0] Accum2_acc_1785_nl;
  wire[16:0] nl_Accum2_acc_1785_nl;
  wire[19:0] Product1_2_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_2_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_3_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_3_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1784_nl;
  wire[16:0] nl_Accum2_acc_1784_nl;
  wire[19:0] Product1_4_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_4_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_5_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_5_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1783_nl;
  wire[16:0] nl_Accum2_acc_1783_nl;
  wire[19:0] Product1_6_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_6_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_7_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_7_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1782_nl;
  wire[16:0] nl_Accum2_acc_1782_nl;
  wire[19:0] Product1_8_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_8_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_9_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_9_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1790_nl;
  wire[16:0] nl_Accum2_acc_1790_nl;
  wire[15:0] Accum2_acc_1787_nl;
  wire[16:0] nl_Accum2_acc_1787_nl;
  wire[15:0] Accum2_acc_1781_nl;
  wire[16:0] nl_Accum2_acc_1781_nl;
  wire[19:0] Product1_10_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_10_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_11_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_11_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1780_nl;
  wire[16:0] nl_Accum2_acc_1780_nl;
  wire[19:0] Product1_12_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_12_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_13_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_13_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[15:0] Accum2_acc_1786_nl;
  wire[16:0] nl_Accum2_acc_1786_nl;
  wire[9:0] Accum2_acc_1919_nl;
  wire[10:0] nl_Accum2_acc_1919_nl;
  wire[19:0] Product1_1_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_1_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[14:0] Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[16:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[19:0] Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[19:0] Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire signed [20:0] nl_Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [47:0] nl_layer6_out_rsci_idat;
  assign nl_layer6_out_rsci_idat = {layer6_out_rsci_idat_47_32 , layer6_out_rsci_idat_31_16
      , layer6_out_rsci_idat_15_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd224)) input_1_rsci (
      .dat(input_1_rsc_dat),
      .idat(input_1_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd48)) layer6_out_rsci (
      .idat(nl_layer6_out_rsci_idat[47:0]),
      .dat(layer6_out_rsc_dat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd8960)) w2_rsci (
      .dat(w2_rsc_dat),
      .idat(w2_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd640)) b2_rsci (
      .dat(b2_rsc_dat),
      .idat(b2_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd1920)) w5_rsci (
      .dat(w5_rsc_dat),
      .idat(w5_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd15)) b5_rsci (
      .dat(b5_rsc_dat),
      .idat(b5_rsci_idat)
    );
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[644:640]));
  assign Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1284:1280]));
  assign Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_134_nl = (readslicef_20_16_4(Product1_2_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_134_nl = nl_Accum2_acc_134_nl[15:0];
  assign nl_Product1_4_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1924:1920]));
  assign Product1_4_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2564:2560]));
  assign Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_133_nl = (readslicef_20_16_4(Product1_4_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_133_nl = nl_Accum2_acc_133_nl[15:0];
  assign nl_Product1_6_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3204:3200]));
  assign Product1_6_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3844:3840]));
  assign Product1_7_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_132_nl = (readslicef_20_16_4(Product1_6_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_132_nl = nl_Accum2_acc_132_nl[15:0];
  assign nl_Product1_8_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4484:4480]));
  assign Product1_8_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5124:5120]));
  assign Product1_9_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_131_nl = (readslicef_20_16_4(Product1_8_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_131_nl = nl_Accum2_acc_131_nl[15:0];
  assign nl_Accum2_acc_140_nl = Accum2_acc_134_nl + Accum2_acc_133_nl + Accum2_acc_132_nl
      + Accum2_acc_131_nl;
  assign Accum2_acc_140_nl = nl_Accum2_acc_140_nl[15:0];
  assign nl_Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5764:5760]));
  assign Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6404:6400]));
  assign Product1_11_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_130_nl = (readslicef_20_16_4(Product1_10_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_130_nl = nl_Accum2_acc_130_nl[15:0];
  assign nl_Product1_12_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7044:7040]));
  assign Product1_12_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7684:7680]));
  assign Product1_13_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_129_nl = (readslicef_20_16_4(Product1_12_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_129_nl = nl_Accum2_acc_129_nl[15:0];
  assign nl_Accum2_acc_136_nl = Accum2_acc_130_nl + Accum2_acc_129_nl;
  assign Accum2_acc_136_nl = nl_Accum2_acc_136_nl[15:0];
  assign nl_Accum2_acc_1792_nl = (Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[4:0]);
  assign Accum2_acc_1792_nl = nl_Accum2_acc_1792_nl[9:0];
  assign nl_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[4:0]));
  assign Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_139_nl = ({Accum2_acc_1792_nl , (Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_139_nl = nl_Accum2_acc_139_nl[15:0];
  assign nl_Accum2_acc_nl = Accum2_acc_136_nl + Accum2_acc_139_nl;
  assign Accum2_acc_nl = nl_Accum2_acc_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1 = Accum2_acc_140_nl
      + Accum2_acc_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[649:645]));
  assign Product1_2_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1289:1285]));
  assign Product1_3_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_147_nl = (readslicef_20_16_4(Product1_2_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_147_nl = nl_Accum2_acc_147_nl[15:0];
  assign nl_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1929:1925]));
  assign Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2569:2565]));
  assign Product1_5_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_146_nl = (readslicef_20_16_4(Product1_4_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_146_nl = nl_Accum2_acc_146_nl[15:0];
  assign nl_Product1_6_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3209:3205]));
  assign Product1_6_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3849:3845]));
  assign Product1_7_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_145_nl = (readslicef_20_16_4(Product1_6_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_145_nl = nl_Accum2_acc_145_nl[15:0];
  assign nl_Product1_8_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4489:4485]));
  assign Product1_8_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5129:5125]));
  assign Product1_9_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_144_nl = (readslicef_20_16_4(Product1_8_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_144_nl = nl_Accum2_acc_144_nl[15:0];
  assign nl_Accum2_acc_153_nl = Accum2_acc_147_nl + Accum2_acc_146_nl + Accum2_acc_145_nl
      + Accum2_acc_144_nl;
  assign Accum2_acc_153_nl = nl_Accum2_acc_153_nl[15:0];
  assign nl_Product1_10_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5769:5765]));
  assign Product1_10_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6409:6405]));
  assign Product1_11_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_143_nl = (readslicef_20_16_4(Product1_10_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_143_nl = nl_Accum2_acc_143_nl[15:0];
  assign nl_Product1_12_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7049:7045]));
  assign Product1_12_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7689:7685]));
  assign Product1_13_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_142_nl = (readslicef_20_16_4(Product1_12_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_142_nl = nl_Accum2_acc_142_nl[15:0];
  assign nl_Accum2_acc_149_nl = Accum2_acc_143_nl + Accum2_acc_142_nl;
  assign Accum2_acc_149_nl = nl_Accum2_acc_149_nl[15:0];
  assign nl_Accum2_acc_1793_nl = (Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[9:5]);
  assign Accum2_acc_1793_nl = nl_Accum2_acc_1793_nl[9:0];
  assign nl_Product1_1_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[9:5]));
  assign Product1_1_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_148_nl = ({Accum2_acc_1793_nl , (Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_148_nl = nl_Accum2_acc_148_nl[15:0];
  assign nl_Accum2_acc_152_nl = Accum2_acc_149_nl + Accum2_acc_148_nl;
  assign Accum2_acc_152_nl = nl_Accum2_acc_152_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1 = Accum2_acc_153_nl
      + Accum2_acc_152_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[654:650]));
  assign Product1_2_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1294:1290]));
  assign Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_160_nl = (readslicef_20_16_4(Product1_2_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_160_nl = nl_Accum2_acc_160_nl[15:0];
  assign nl_Product1_4_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1934:1930]));
  assign Product1_4_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2574:2570]));
  assign Product1_5_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_159_nl = (readslicef_20_16_4(Product1_4_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_159_nl = nl_Accum2_acc_159_nl[15:0];
  assign nl_Product1_6_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3214:3210]));
  assign Product1_6_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3854:3850]));
  assign Product1_7_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_158_nl = (readslicef_20_16_4(Product1_6_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_158_nl = nl_Accum2_acc_158_nl[15:0];
  assign nl_Product1_8_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4494:4490]));
  assign Product1_8_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5134:5130]));
  assign Product1_9_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_157_nl = (readslicef_20_16_4(Product1_8_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_157_nl = nl_Accum2_acc_157_nl[15:0];
  assign nl_Accum2_acc_166_nl = Accum2_acc_160_nl + Accum2_acc_159_nl + Accum2_acc_158_nl
      + Accum2_acc_157_nl;
  assign Accum2_acc_166_nl = nl_Accum2_acc_166_nl[15:0];
  assign nl_Product1_10_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5774:5770]));
  assign Product1_10_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6414:6410]));
  assign Product1_11_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_156_nl = (readslicef_20_16_4(Product1_10_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_156_nl = nl_Accum2_acc_156_nl[15:0];
  assign nl_Product1_12_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7054:7050]));
  assign Product1_12_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7694:7690]));
  assign Product1_13_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_155_nl = (readslicef_20_16_4(Product1_12_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_155_nl = nl_Accum2_acc_155_nl[15:0];
  assign nl_Accum2_acc_162_nl = Accum2_acc_156_nl + Accum2_acc_155_nl;
  assign Accum2_acc_162_nl = nl_Accum2_acc_162_nl[15:0];
  assign nl_Accum2_acc_1794_nl = (Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[14:10]);
  assign Accum2_acc_1794_nl = nl_Accum2_acc_1794_nl[9:0];
  assign nl_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[14:10]));
  assign Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_161_nl = ({Accum2_acc_1794_nl , (Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_161_nl = nl_Accum2_acc_161_nl[15:0];
  assign nl_Accum2_acc_165_nl = Accum2_acc_162_nl + Accum2_acc_161_nl;
  assign Accum2_acc_165_nl = nl_Accum2_acc_165_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1 = Accum2_acc_166_nl
      + Accum2_acc_165_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[659:655]));
  assign Product1_2_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1299:1295]));
  assign Product1_3_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_173_nl = (readslicef_20_16_4(Product1_2_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_173_nl = nl_Accum2_acc_173_nl[15:0];
  assign nl_Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1939:1935]));
  assign Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2579:2575]));
  assign Product1_5_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_172_nl = (readslicef_20_16_4(Product1_4_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_172_nl = nl_Accum2_acc_172_nl[15:0];
  assign nl_Product1_6_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3219:3215]));
  assign Product1_6_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3859:3855]));
  assign Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_171_nl = (readslicef_20_16_4(Product1_6_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_171_nl = nl_Accum2_acc_171_nl[15:0];
  assign nl_Product1_8_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4499:4495]));
  assign Product1_8_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5139:5135]));
  assign Product1_9_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_170_nl = (readslicef_20_16_4(Product1_8_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_170_nl = nl_Accum2_acc_170_nl[15:0];
  assign nl_Accum2_acc_179_nl = Accum2_acc_173_nl + Accum2_acc_172_nl + Accum2_acc_171_nl
      + Accum2_acc_170_nl;
  assign Accum2_acc_179_nl = nl_Accum2_acc_179_nl[15:0];
  assign nl_Product1_10_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5779:5775]));
  assign Product1_10_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6419:6415]));
  assign Product1_11_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_169_nl = (readslicef_20_16_4(Product1_10_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_169_nl = nl_Accum2_acc_169_nl[15:0];
  assign nl_Product1_12_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7059:7055]));
  assign Product1_12_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7699:7695]));
  assign Product1_13_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_168_nl = (readslicef_20_16_4(Product1_12_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_168_nl = nl_Accum2_acc_168_nl[15:0];
  assign nl_Accum2_acc_175_nl = Accum2_acc_169_nl + Accum2_acc_168_nl;
  assign Accum2_acc_175_nl = nl_Accum2_acc_175_nl[15:0];
  assign nl_Accum2_acc_1795_nl = (Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[19:15]);
  assign Accum2_acc_1795_nl = nl_Accum2_acc_1795_nl[9:0];
  assign nl_Product1_1_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[19:15]));
  assign Product1_1_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_174_nl = ({Accum2_acc_1795_nl , (Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_174_nl = nl_Accum2_acc_174_nl[15:0];
  assign nl_Accum2_acc_178_nl = Accum2_acc_175_nl + Accum2_acc_174_nl;
  assign Accum2_acc_178_nl = nl_Accum2_acc_178_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1 = Accum2_acc_179_nl
      + Accum2_acc_178_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[664:660]));
  assign Product1_2_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1304:1300]));
  assign Product1_3_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_186_nl = (readslicef_20_16_4(Product1_2_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_186_nl = nl_Accum2_acc_186_nl[15:0];
  assign nl_Product1_4_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1944:1940]));
  assign Product1_4_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2584:2580]));
  assign Product1_5_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_185_nl = (readslicef_20_16_4(Product1_4_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_185_nl = nl_Accum2_acc_185_nl[15:0];
  assign nl_Product1_6_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3224:3220]));
  assign Product1_6_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3864:3860]));
  assign Product1_7_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_184_nl = (readslicef_20_16_4(Product1_6_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_184_nl = nl_Accum2_acc_184_nl[15:0];
  assign nl_Product1_8_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4504:4500]));
  assign Product1_8_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5144:5140]));
  assign Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_183_nl = (readslicef_20_16_4(Product1_8_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_183_nl = nl_Accum2_acc_183_nl[15:0];
  assign nl_Accum2_acc_192_nl = Accum2_acc_186_nl + Accum2_acc_185_nl + Accum2_acc_184_nl
      + Accum2_acc_183_nl;
  assign Accum2_acc_192_nl = nl_Accum2_acc_192_nl[15:0];
  assign nl_Product1_10_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5784:5780]));
  assign Product1_10_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6424:6420]));
  assign Product1_11_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_182_nl = (readslicef_20_16_4(Product1_10_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_182_nl = nl_Accum2_acc_182_nl[15:0];
  assign nl_Product1_12_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7064:7060]));
  assign Product1_12_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7704:7700]));
  assign Product1_13_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_181_nl = (readslicef_20_16_4(Product1_12_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_181_nl = nl_Accum2_acc_181_nl[15:0];
  assign nl_Accum2_acc_188_nl = Accum2_acc_182_nl + Accum2_acc_181_nl;
  assign Accum2_acc_188_nl = nl_Accum2_acc_188_nl[15:0];
  assign nl_Accum2_acc_1796_nl = (Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[24:20]);
  assign Accum2_acc_1796_nl = nl_Accum2_acc_1796_nl[9:0];
  assign nl_Product1_1_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[24:20]));
  assign Product1_1_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_187_nl = ({Accum2_acc_1796_nl , (Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_187_nl = nl_Accum2_acc_187_nl[15:0];
  assign nl_Accum2_acc_191_nl = Accum2_acc_188_nl + Accum2_acc_187_nl;
  assign Accum2_acc_191_nl = nl_Accum2_acc_191_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1 = Accum2_acc_192_nl
      + Accum2_acc_191_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[669:665]));
  assign Product1_2_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1309:1305]));
  assign Product1_3_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_199_nl = (readslicef_20_16_4(Product1_2_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_199_nl = nl_Accum2_acc_199_nl[15:0];
  assign nl_Product1_4_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1949:1945]));
  assign Product1_4_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2589:2585]));
  assign Product1_5_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_198_nl = (readslicef_20_16_4(Product1_4_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_198_nl = nl_Accum2_acc_198_nl[15:0];
  assign nl_Product1_6_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3229:3225]));
  assign Product1_6_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3869:3865]));
  assign Product1_7_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_197_nl = (readslicef_20_16_4(Product1_6_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_197_nl = nl_Accum2_acc_197_nl[15:0];
  assign nl_Product1_8_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4509:4505]));
  assign Product1_8_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5149:5145]));
  assign Product1_9_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_196_nl = (readslicef_20_16_4(Product1_8_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_196_nl = nl_Accum2_acc_196_nl[15:0];
  assign nl_Accum2_acc_205_nl = Accum2_acc_199_nl + Accum2_acc_198_nl + Accum2_acc_197_nl
      + Accum2_acc_196_nl;
  assign Accum2_acc_205_nl = nl_Accum2_acc_205_nl[15:0];
  assign nl_Product1_10_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5789:5785]));
  assign Product1_10_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6429:6425]));
  assign Product1_11_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_195_nl = (readslicef_20_16_4(Product1_10_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_195_nl = nl_Accum2_acc_195_nl[15:0];
  assign nl_Product1_12_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7069:7065]));
  assign Product1_12_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7709:7705]));
  assign Product1_13_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_194_nl = (readslicef_20_16_4(Product1_12_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_194_nl = nl_Accum2_acc_194_nl[15:0];
  assign nl_Accum2_acc_201_nl = Accum2_acc_195_nl + Accum2_acc_194_nl;
  assign Accum2_acc_201_nl = nl_Accum2_acc_201_nl[15:0];
  assign nl_Accum2_acc_1797_nl = (Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[29:25]);
  assign Accum2_acc_1797_nl = nl_Accum2_acc_1797_nl[9:0];
  assign nl_Product1_1_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[29:25]));
  assign Product1_1_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_200_nl = ({Accum2_acc_1797_nl , (Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_200_nl = nl_Accum2_acc_200_nl[15:0];
  assign nl_Accum2_acc_204_nl = Accum2_acc_201_nl + Accum2_acc_200_nl;
  assign Accum2_acc_204_nl = nl_Accum2_acc_204_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1 = Accum2_acc_205_nl
      + Accum2_acc_204_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[674:670]));
  assign Product1_2_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1314:1310]));
  assign Product1_3_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_212_nl = (readslicef_20_16_4(Product1_2_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_212_nl = nl_Accum2_acc_212_nl[15:0];
  assign nl_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1954:1950]));
  assign Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2594:2590]));
  assign Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_211_nl = (readslicef_20_16_4(Product1_4_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_211_nl = nl_Accum2_acc_211_nl[15:0];
  assign nl_Product1_6_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3234:3230]));
  assign Product1_6_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3874:3870]));
  assign Product1_7_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_210_nl = (readslicef_20_16_4(Product1_6_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_210_nl = nl_Accum2_acc_210_nl[15:0];
  assign nl_Product1_8_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4514:4510]));
  assign Product1_8_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5154:5150]));
  assign Product1_9_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_209_nl = (readslicef_20_16_4(Product1_8_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_209_nl = nl_Accum2_acc_209_nl[15:0];
  assign nl_Accum2_acc_218_nl = Accum2_acc_212_nl + Accum2_acc_211_nl + Accum2_acc_210_nl
      + Accum2_acc_209_nl;
  assign Accum2_acc_218_nl = nl_Accum2_acc_218_nl[15:0];
  assign nl_Product1_10_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5794:5790]));
  assign Product1_10_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6434:6430]));
  assign Product1_11_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_208_nl = (readslicef_20_16_4(Product1_10_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_208_nl = nl_Accum2_acc_208_nl[15:0];
  assign nl_Product1_12_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7074:7070]));
  assign Product1_12_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7714:7710]));
  assign Product1_13_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_207_nl = (readslicef_20_16_4(Product1_12_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_207_nl = nl_Accum2_acc_207_nl[15:0];
  assign nl_Accum2_acc_214_nl = Accum2_acc_208_nl + Accum2_acc_207_nl;
  assign Accum2_acc_214_nl = nl_Accum2_acc_214_nl[15:0];
  assign nl_Accum2_acc_1798_nl = (Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[34:30]);
  assign Accum2_acc_1798_nl = nl_Accum2_acc_1798_nl[9:0];
  assign nl_Product1_1_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[34:30]));
  assign Product1_1_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_213_nl = ({Accum2_acc_1798_nl , (Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_213_nl = nl_Accum2_acc_213_nl[15:0];
  assign nl_Accum2_acc_217_nl = Accum2_acc_214_nl + Accum2_acc_213_nl;
  assign Accum2_acc_217_nl = nl_Accum2_acc_217_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1 = Accum2_acc_218_nl
      + Accum2_acc_217_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[679:675]));
  assign Product1_2_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1319:1315]));
  assign Product1_3_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_225_nl = (readslicef_20_16_4(Product1_2_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_225_nl = nl_Accum2_acc_225_nl[15:0];
  assign nl_Product1_4_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1959:1955]));
  assign Product1_4_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2599:2595]));
  assign Product1_5_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_224_nl = (readslicef_20_16_4(Product1_4_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_224_nl = nl_Accum2_acc_224_nl[15:0];
  assign nl_Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3239:3235]));
  assign Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3879:3875]));
  assign Product1_7_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_223_nl = (readslicef_20_16_4(Product1_6_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_223_nl = nl_Accum2_acc_223_nl[15:0];
  assign nl_Product1_8_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4519:4515]));
  assign Product1_8_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5159:5155]));
  assign Product1_9_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_222_nl = (readslicef_20_16_4(Product1_8_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_222_nl = nl_Accum2_acc_222_nl[15:0];
  assign nl_Accum2_acc_231_nl = Accum2_acc_225_nl + Accum2_acc_224_nl + Accum2_acc_223_nl
      + Accum2_acc_222_nl;
  assign Accum2_acc_231_nl = nl_Accum2_acc_231_nl[15:0];
  assign nl_Product1_10_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5799:5795]));
  assign Product1_10_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6439:6435]));
  assign Product1_11_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_221_nl = (readslicef_20_16_4(Product1_10_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_221_nl = nl_Accum2_acc_221_nl[15:0];
  assign nl_Product1_12_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7079:7075]));
  assign Product1_12_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7719:7715]));
  assign Product1_13_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_220_nl = (readslicef_20_16_4(Product1_12_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_220_nl = nl_Accum2_acc_220_nl[15:0];
  assign nl_Accum2_acc_227_nl = Accum2_acc_221_nl + Accum2_acc_220_nl;
  assign Accum2_acc_227_nl = nl_Accum2_acc_227_nl[15:0];
  assign nl_Accum2_acc_1799_nl = (Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[39:35]);
  assign Accum2_acc_1799_nl = nl_Accum2_acc_1799_nl[9:0];
  assign nl_Product1_1_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[39:35]));
  assign Product1_1_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_226_nl = ({Accum2_acc_1799_nl , (Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_226_nl = nl_Accum2_acc_226_nl[15:0];
  assign nl_Accum2_acc_230_nl = Accum2_acc_227_nl + Accum2_acc_226_nl;
  assign Accum2_acc_230_nl = nl_Accum2_acc_230_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1 = Accum2_acc_231_nl
      + Accum2_acc_230_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[684:680]));
  assign Product1_2_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1324:1320]));
  assign Product1_3_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_238_nl = (readslicef_20_16_4(Product1_2_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_238_nl = nl_Accum2_acc_238_nl[15:0];
  assign nl_Product1_4_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1964:1960]));
  assign Product1_4_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2604:2600]));
  assign Product1_5_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_237_nl = (readslicef_20_16_4(Product1_4_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_237_nl = nl_Accum2_acc_237_nl[15:0];
  assign nl_Product1_6_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3244:3240]));
  assign Product1_6_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3884:3880]));
  assign Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_236_nl = (readslicef_20_16_4(Product1_6_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_236_nl = nl_Accum2_acc_236_nl[15:0];
  assign nl_Product1_8_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4524:4520]));
  assign Product1_8_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5164:5160]));
  assign Product1_9_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_235_nl = (readslicef_20_16_4(Product1_8_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_235_nl = nl_Accum2_acc_235_nl[15:0];
  assign nl_Accum2_acc_244_nl = Accum2_acc_238_nl + Accum2_acc_237_nl + Accum2_acc_236_nl
      + Accum2_acc_235_nl;
  assign Accum2_acc_244_nl = nl_Accum2_acc_244_nl[15:0];
  assign nl_Product1_10_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5804:5800]));
  assign Product1_10_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6444:6440]));
  assign Product1_11_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_234_nl = (readslicef_20_16_4(Product1_10_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_234_nl = nl_Accum2_acc_234_nl[15:0];
  assign nl_Product1_12_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7084:7080]));
  assign Product1_12_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7724:7720]));
  assign Product1_13_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_233_nl = (readslicef_20_16_4(Product1_12_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_233_nl = nl_Accum2_acc_233_nl[15:0];
  assign nl_Accum2_acc_240_nl = Accum2_acc_234_nl + Accum2_acc_233_nl;
  assign Accum2_acc_240_nl = nl_Accum2_acc_240_nl[15:0];
  assign nl_Accum2_acc_1800_nl = (Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[44:40]);
  assign Accum2_acc_1800_nl = nl_Accum2_acc_1800_nl[9:0];
  assign nl_Product1_1_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[44:40]));
  assign Product1_1_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_239_nl = ({Accum2_acc_1800_nl , (Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_239_nl = nl_Accum2_acc_239_nl[15:0];
  assign nl_Accum2_acc_243_nl = Accum2_acc_240_nl + Accum2_acc_239_nl;
  assign Accum2_acc_243_nl = nl_Accum2_acc_243_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1 = Accum2_acc_244_nl
      + Accum2_acc_243_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[689:685]));
  assign Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1329:1325]));
  assign Product1_3_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_251_nl = (readslicef_20_16_4(Product1_2_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_251_nl = nl_Accum2_acc_251_nl[15:0];
  assign nl_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1969:1965]));
  assign Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2609:2605]));
  assign Product1_5_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_250_nl = (readslicef_20_16_4(Product1_4_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_250_nl = nl_Accum2_acc_250_nl[15:0];
  assign nl_Product1_6_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3249:3245]));
  assign Product1_6_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3889:3885]));
  assign Product1_7_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_249_nl = (readslicef_20_16_4(Product1_6_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_249_nl = nl_Accum2_acc_249_nl[15:0];
  assign nl_Product1_8_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4529:4525]));
  assign Product1_8_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5169:5165]));
  assign Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_248_nl = (readslicef_20_16_4(Product1_8_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_248_nl = nl_Accum2_acc_248_nl[15:0];
  assign nl_Accum2_acc_257_nl = Accum2_acc_251_nl + Accum2_acc_250_nl + Accum2_acc_249_nl
      + Accum2_acc_248_nl;
  assign Accum2_acc_257_nl = nl_Accum2_acc_257_nl[15:0];
  assign nl_Product1_10_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5809:5805]));
  assign Product1_10_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6449:6445]));
  assign Product1_11_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_247_nl = (readslicef_20_16_4(Product1_10_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_247_nl = nl_Accum2_acc_247_nl[15:0];
  assign nl_Product1_12_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7089:7085]));
  assign Product1_12_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7729:7725]));
  assign Product1_13_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_246_nl = (readslicef_20_16_4(Product1_12_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_246_nl = nl_Accum2_acc_246_nl[15:0];
  assign nl_Accum2_acc_253_nl = Accum2_acc_247_nl + Accum2_acc_246_nl;
  assign Accum2_acc_253_nl = nl_Accum2_acc_253_nl[15:0];
  assign nl_Accum2_acc_1801_nl = (Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[49:45]);
  assign Accum2_acc_1801_nl = nl_Accum2_acc_1801_nl[9:0];
  assign nl_Product1_1_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[49:45]));
  assign Product1_1_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_252_nl = ({Accum2_acc_1801_nl , (Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_252_nl = nl_Accum2_acc_252_nl[15:0];
  assign nl_Accum2_acc_256_nl = Accum2_acc_253_nl + Accum2_acc_252_nl;
  assign Accum2_acc_256_nl = nl_Accum2_acc_256_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1 = Accum2_acc_257_nl
      + Accum2_acc_256_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[694:690]));
  assign Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1334:1330]));
  assign Product1_3_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_264_nl = (readslicef_20_16_4(Product1_2_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_264_nl = nl_Accum2_acc_264_nl[15:0];
  assign nl_Product1_4_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1974:1970]));
  assign Product1_4_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2614:2610]));
  assign Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_263_nl = (readslicef_20_16_4(Product1_4_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_263_nl = nl_Accum2_acc_263_nl[15:0];
  assign nl_Product1_6_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3254:3250]));
  assign Product1_6_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3894:3890]));
  assign Product1_7_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_262_nl = (readslicef_20_16_4(Product1_6_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_262_nl = nl_Accum2_acc_262_nl[15:0];
  assign nl_Product1_8_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4534:4530]));
  assign Product1_8_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5174:5170]));
  assign Product1_9_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_261_nl = (readslicef_20_16_4(Product1_8_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_261_nl = nl_Accum2_acc_261_nl[15:0];
  assign nl_Accum2_acc_270_nl = Accum2_acc_264_nl + Accum2_acc_263_nl + Accum2_acc_262_nl
      + Accum2_acc_261_nl;
  assign Accum2_acc_270_nl = nl_Accum2_acc_270_nl[15:0];
  assign nl_Product1_10_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5814:5810]));
  assign Product1_10_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6454:6450]));
  assign Product1_11_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_260_nl = (readslicef_20_16_4(Product1_10_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_260_nl = nl_Accum2_acc_260_nl[15:0];
  assign nl_Product1_12_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7094:7090]));
  assign Product1_12_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7734:7730]));
  assign Product1_13_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_259_nl = (readslicef_20_16_4(Product1_12_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_259_nl = nl_Accum2_acc_259_nl[15:0];
  assign nl_Accum2_acc_266_nl = Accum2_acc_260_nl + Accum2_acc_259_nl;
  assign Accum2_acc_266_nl = nl_Accum2_acc_266_nl[15:0];
  assign nl_Accum2_acc_1802_nl = (Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[54:50]);
  assign Accum2_acc_1802_nl = nl_Accum2_acc_1802_nl[9:0];
  assign nl_Product1_1_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[54:50]));
  assign Product1_1_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_265_nl = ({Accum2_acc_1802_nl , (Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_265_nl = nl_Accum2_acc_265_nl[15:0];
  assign nl_Accum2_acc_269_nl = Accum2_acc_266_nl + Accum2_acc_265_nl;
  assign Accum2_acc_269_nl = nl_Accum2_acc_269_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1 = Accum2_acc_270_nl
      + Accum2_acc_269_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[699:695]));
  assign Product1_2_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1339:1335]));
  assign Product1_3_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_277_nl = (readslicef_20_16_4(Product1_2_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_277_nl = nl_Accum2_acc_277_nl[15:0];
  assign nl_Product1_4_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1979:1975]));
  assign Product1_4_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2619:2615]));
  assign Product1_5_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_276_nl = (readslicef_20_16_4(Product1_4_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_276_nl = nl_Accum2_acc_276_nl[15:0];
  assign nl_Product1_6_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3259:3255]));
  assign Product1_6_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3899:3895]));
  assign Product1_7_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_275_nl = (readslicef_20_16_4(Product1_6_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_275_nl = nl_Accum2_acc_275_nl[15:0];
  assign nl_Product1_8_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4539:4535]));
  assign Product1_8_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5179:5175]));
  assign Product1_9_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_274_nl = (readslicef_20_16_4(Product1_8_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_274_nl = nl_Accum2_acc_274_nl[15:0];
  assign nl_Accum2_acc_283_nl = Accum2_acc_277_nl + Accum2_acc_276_nl + Accum2_acc_275_nl
      + Accum2_acc_274_nl;
  assign Accum2_acc_283_nl = nl_Accum2_acc_283_nl[15:0];
  assign nl_Product1_10_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5819:5815]));
  assign Product1_10_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6459:6455]));
  assign Product1_11_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_273_nl = (readslicef_20_16_4(Product1_10_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_273_nl = nl_Accum2_acc_273_nl[15:0];
  assign nl_Product1_12_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7099:7095]));
  assign Product1_12_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7739:7735]));
  assign Product1_13_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_272_nl = (readslicef_20_16_4(Product1_12_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_272_nl = nl_Accum2_acc_272_nl[15:0];
  assign nl_Accum2_acc_279_nl = Accum2_acc_273_nl + Accum2_acc_272_nl;
  assign Accum2_acc_279_nl = nl_Accum2_acc_279_nl[15:0];
  assign nl_Accum2_acc_1803_nl = (Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[59:55]);
  assign Accum2_acc_1803_nl = nl_Accum2_acc_1803_nl[9:0];
  assign nl_Product1_1_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[59:55]));
  assign Product1_1_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_278_nl = ({Accum2_acc_1803_nl , (Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_278_nl = nl_Accum2_acc_278_nl[15:0];
  assign nl_Accum2_acc_282_nl = Accum2_acc_279_nl + Accum2_acc_278_nl;
  assign Accum2_acc_282_nl = nl_Accum2_acc_282_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1 = Accum2_acc_283_nl
      + Accum2_acc_282_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[704:700]));
  assign Product1_2_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1344:1340]));
  assign Product1_3_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_290_nl = (readslicef_20_16_4(Product1_2_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_290_nl = nl_Accum2_acc_290_nl[15:0];
  assign nl_Product1_4_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1984:1980]));
  assign Product1_4_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2624:2620]));
  assign Product1_5_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_289_nl = (readslicef_20_16_4(Product1_4_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_289_nl = nl_Accum2_acc_289_nl[15:0];
  assign nl_Product1_6_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3264:3260]));
  assign Product1_6_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3904:3900]));
  assign Product1_7_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_288_nl = (readslicef_20_16_4(Product1_6_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_288_nl = nl_Accum2_acc_288_nl[15:0];
  assign nl_Product1_8_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4544:4540]));
  assign Product1_8_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5184:5180]));
  assign Product1_9_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_287_nl = (readslicef_20_16_4(Product1_8_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_287_nl = nl_Accum2_acc_287_nl[15:0];
  assign nl_Accum2_acc_296_nl = Accum2_acc_290_nl + Accum2_acc_289_nl + Accum2_acc_288_nl
      + Accum2_acc_287_nl;
  assign Accum2_acc_296_nl = nl_Accum2_acc_296_nl[15:0];
  assign nl_Product1_10_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5824:5820]));
  assign Product1_10_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6464:6460]));
  assign Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_286_nl = (readslicef_20_16_4(Product1_10_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_286_nl = nl_Accum2_acc_286_nl[15:0];
  assign nl_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7104:7100]));
  assign Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7744:7740]));
  assign Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_285_nl = (readslicef_20_16_4(Product1_12_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_285_nl = nl_Accum2_acc_285_nl[15:0];
  assign nl_Accum2_acc_292_nl = Accum2_acc_286_nl + Accum2_acc_285_nl;
  assign Accum2_acc_292_nl = nl_Accum2_acc_292_nl[15:0];
  assign nl_Accum2_acc_1804_nl = (Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[64:60]);
  assign Accum2_acc_1804_nl = nl_Accum2_acc_1804_nl[9:0];
  assign nl_Product1_1_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[64:60]));
  assign Product1_1_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_291_nl = ({Accum2_acc_1804_nl , (Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_291_nl = nl_Accum2_acc_291_nl[15:0];
  assign nl_Accum2_acc_295_nl = Accum2_acc_292_nl + Accum2_acc_291_nl;
  assign Accum2_acc_295_nl = nl_Accum2_acc_295_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1 = Accum2_acc_296_nl
      + Accum2_acc_295_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[709:705]));
  assign Product1_2_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1349:1345]));
  assign Product1_3_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_303_nl = (readslicef_20_16_4(Product1_2_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_303_nl = nl_Accum2_acc_303_nl[15:0];
  assign nl_Product1_4_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1989:1985]));
  assign Product1_4_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2629:2625]));
  assign Product1_5_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_302_nl = (readslicef_20_16_4(Product1_4_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_302_nl = nl_Accum2_acc_302_nl[15:0];
  assign nl_Product1_6_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3269:3265]));
  assign Product1_6_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3909:3905]));
  assign Product1_7_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_301_nl = (readslicef_20_16_4(Product1_6_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_301_nl = nl_Accum2_acc_301_nl[15:0];
  assign nl_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4549:4545]));
  assign Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5189:5185]));
  assign Product1_9_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_300_nl = (readslicef_20_16_4(Product1_8_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_300_nl = nl_Accum2_acc_300_nl[15:0];
  assign nl_Accum2_acc_309_nl = Accum2_acc_303_nl + Accum2_acc_302_nl + Accum2_acc_301_nl
      + Accum2_acc_300_nl;
  assign Accum2_acc_309_nl = nl_Accum2_acc_309_nl[15:0];
  assign nl_Product1_10_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5829:5825]));
  assign Product1_10_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6469:6465]));
  assign Product1_11_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_299_nl = (readslicef_20_16_4(Product1_10_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_299_nl = nl_Accum2_acc_299_nl[15:0];
  assign nl_Product1_12_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7109:7105]));
  assign Product1_12_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7749:7745]));
  assign Product1_13_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_298_nl = (readslicef_20_16_4(Product1_12_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_298_nl = nl_Accum2_acc_298_nl[15:0];
  assign nl_Accum2_acc_305_nl = Accum2_acc_299_nl + Accum2_acc_298_nl;
  assign Accum2_acc_305_nl = nl_Accum2_acc_305_nl[15:0];
  assign nl_Accum2_acc_1805_nl = (Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[69:65]);
  assign Accum2_acc_1805_nl = nl_Accum2_acc_1805_nl[9:0];
  assign nl_Product1_1_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[69:65]));
  assign Product1_1_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_304_nl = ({Accum2_acc_1805_nl , (Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_304_nl = nl_Accum2_acc_304_nl[15:0];
  assign nl_Accum2_acc_308_nl = Accum2_acc_305_nl + Accum2_acc_304_nl;
  assign Accum2_acc_308_nl = nl_Accum2_acc_308_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1 = Accum2_acc_309_nl
      + Accum2_acc_308_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[714:710]));
  assign Product1_2_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1354:1350]));
  assign Product1_3_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_316_nl = (readslicef_20_16_4(Product1_2_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_316_nl = nl_Accum2_acc_316_nl[15:0];
  assign nl_Product1_4_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1994:1990]));
  assign Product1_4_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2634:2630]));
  assign Product1_5_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_315_nl = (readslicef_20_16_4(Product1_4_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_315_nl = nl_Accum2_acc_315_nl[15:0];
  assign nl_Product1_6_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3274:3270]));
  assign Product1_6_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3914:3910]));
  assign Product1_7_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_314_nl = (readslicef_20_16_4(Product1_6_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_314_nl = nl_Accum2_acc_314_nl[15:0];
  assign nl_Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4554:4550]));
  assign Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5194:5190]));
  assign Product1_9_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_313_nl = (readslicef_20_16_4(Product1_8_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_313_nl = nl_Accum2_acc_313_nl[15:0];
  assign nl_Accum2_acc_322_nl = Accum2_acc_316_nl + Accum2_acc_315_nl + Accum2_acc_314_nl
      + Accum2_acc_313_nl;
  assign Accum2_acc_322_nl = nl_Accum2_acc_322_nl[15:0];
  assign nl_Product1_10_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5834:5830]));
  assign Product1_10_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6474:6470]));
  assign Product1_11_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_312_nl = (readslicef_20_16_4(Product1_10_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_312_nl = nl_Accum2_acc_312_nl[15:0];
  assign nl_Product1_12_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7114:7110]));
  assign Product1_12_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7754:7750]));
  assign Product1_13_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_311_nl = (readslicef_20_16_4(Product1_12_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_311_nl = nl_Accum2_acc_311_nl[15:0];
  assign nl_Accum2_acc_318_nl = Accum2_acc_312_nl + Accum2_acc_311_nl;
  assign Accum2_acc_318_nl = nl_Accum2_acc_318_nl[15:0];
  assign nl_Accum2_acc_1806_nl = (Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[74:70]);
  assign Accum2_acc_1806_nl = nl_Accum2_acc_1806_nl[9:0];
  assign nl_Product1_1_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[74:70]));
  assign Product1_1_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_317_nl = ({Accum2_acc_1806_nl , (Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_317_nl = nl_Accum2_acc_317_nl[15:0];
  assign nl_Accum2_acc_321_nl = Accum2_acc_318_nl + Accum2_acc_317_nl;
  assign Accum2_acc_321_nl = nl_Accum2_acc_321_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1 = Accum2_acc_322_nl
      + Accum2_acc_321_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[719:715]));
  assign Product1_2_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1359:1355]));
  assign Product1_3_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_329_nl = (readslicef_20_16_4(Product1_2_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_329_nl = nl_Accum2_acc_329_nl[15:0];
  assign nl_Product1_4_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[1999:1995]));
  assign Product1_4_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2639:2635]));
  assign Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_328_nl = (readslicef_20_16_4(Product1_4_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_328_nl = nl_Accum2_acc_328_nl[15:0];
  assign nl_Product1_6_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3279:3275]));
  assign Product1_6_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3919:3915]));
  assign Product1_7_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_327_nl = (readslicef_20_16_4(Product1_6_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_327_nl = nl_Accum2_acc_327_nl[15:0];
  assign nl_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4559:4555]));
  assign Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5199:5195]));
  assign Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_326_nl = (readslicef_20_16_4(Product1_8_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_326_nl = nl_Accum2_acc_326_nl[15:0];
  assign nl_Accum2_acc_335_nl = Accum2_acc_329_nl + Accum2_acc_328_nl + Accum2_acc_327_nl
      + Accum2_acc_326_nl;
  assign Accum2_acc_335_nl = nl_Accum2_acc_335_nl[15:0];
  assign nl_Product1_10_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5839:5835]));
  assign Product1_10_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6479:6475]));
  assign Product1_11_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_325_nl = (readslicef_20_16_4(Product1_10_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_325_nl = nl_Accum2_acc_325_nl[15:0];
  assign nl_Product1_12_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7119:7115]));
  assign Product1_12_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7759:7755]));
  assign Product1_13_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_324_nl = (readslicef_20_16_4(Product1_12_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_324_nl = nl_Accum2_acc_324_nl[15:0];
  assign nl_Accum2_acc_331_nl = Accum2_acc_325_nl + Accum2_acc_324_nl;
  assign Accum2_acc_331_nl = nl_Accum2_acc_331_nl[15:0];
  assign nl_Accum2_acc_1807_nl = (Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[79:75]);
  assign Accum2_acc_1807_nl = nl_Accum2_acc_1807_nl[9:0];
  assign nl_Product1_1_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[79:75]));
  assign Product1_1_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_330_nl = ({Accum2_acc_1807_nl , (Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_330_nl = nl_Accum2_acc_330_nl[15:0];
  assign nl_Accum2_acc_334_nl = Accum2_acc_331_nl + Accum2_acc_330_nl;
  assign Accum2_acc_334_nl = nl_Accum2_acc_334_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1 = Accum2_acc_335_nl
      + Accum2_acc_334_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[724:720]));
  assign Product1_2_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1364:1360]));
  assign Product1_3_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_342_nl = (readslicef_20_16_4(Product1_2_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_342_nl = nl_Accum2_acc_342_nl[15:0];
  assign nl_Product1_4_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2004:2000]));
  assign Product1_4_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2644:2640]));
  assign Product1_5_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_341_nl = (readslicef_20_16_4(Product1_4_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_341_nl = nl_Accum2_acc_341_nl[15:0];
  assign nl_Product1_6_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3284:3280]));
  assign Product1_6_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3924:3920]));
  assign Product1_7_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_340_nl = (readslicef_20_16_4(Product1_6_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_340_nl = nl_Accum2_acc_340_nl[15:0];
  assign nl_Product1_8_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4564:4560]));
  assign Product1_8_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5204:5200]));
  assign Product1_9_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_339_nl = (readslicef_20_16_4(Product1_8_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_339_nl = nl_Accum2_acc_339_nl[15:0];
  assign nl_Accum2_acc_348_nl = Accum2_acc_342_nl + Accum2_acc_341_nl + Accum2_acc_340_nl
      + Accum2_acc_339_nl;
  assign Accum2_acc_348_nl = nl_Accum2_acc_348_nl[15:0];
  assign nl_Product1_10_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5844:5840]));
  assign Product1_10_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6484:6480]));
  assign Product1_11_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_338_nl = (readslicef_20_16_4(Product1_10_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_338_nl = nl_Accum2_acc_338_nl[15:0];
  assign nl_Product1_12_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7124:7120]));
  assign Product1_12_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7764:7760]));
  assign Product1_13_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_337_nl = (readslicef_20_16_4(Product1_12_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_337_nl = nl_Accum2_acc_337_nl[15:0];
  assign nl_Accum2_acc_344_nl = Accum2_acc_338_nl + Accum2_acc_337_nl;
  assign Accum2_acc_344_nl = nl_Accum2_acc_344_nl[15:0];
  assign nl_Accum2_acc_1808_nl = (Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[84:80]);
  assign Accum2_acc_1808_nl = nl_Accum2_acc_1808_nl[9:0];
  assign nl_Product1_1_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[84:80]));
  assign Product1_1_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_343_nl = ({Accum2_acc_1808_nl , (Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_343_nl = nl_Accum2_acc_343_nl[15:0];
  assign nl_Accum2_acc_347_nl = Accum2_acc_344_nl + Accum2_acc_343_nl;
  assign Accum2_acc_347_nl = nl_Accum2_acc_347_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1 = Accum2_acc_348_nl
      + Accum2_acc_347_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[729:725]));
  assign Product1_2_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1369:1365]));
  assign Product1_3_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_355_nl = (readslicef_20_16_4(Product1_2_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_355_nl = nl_Accum2_acc_355_nl[15:0];
  assign nl_Product1_4_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2009:2005]));
  assign Product1_4_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2649:2645]));
  assign Product1_5_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_354_nl = (readslicef_20_16_4(Product1_4_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_354_nl = nl_Accum2_acc_354_nl[15:0];
  assign nl_Product1_6_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3289:3285]));
  assign Product1_6_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3929:3925]));
  assign Product1_7_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_353_nl = (readslicef_20_16_4(Product1_6_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_353_nl = nl_Accum2_acc_353_nl[15:0];
  assign nl_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4569:4565]));
  assign Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5209:5205]));
  assign Product1_9_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_352_nl = (readslicef_20_16_4(Product1_8_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_352_nl = nl_Accum2_acc_352_nl[15:0];
  assign nl_Accum2_acc_361_nl = Accum2_acc_355_nl + Accum2_acc_354_nl + Accum2_acc_353_nl
      + Accum2_acc_352_nl;
  assign Accum2_acc_361_nl = nl_Accum2_acc_361_nl[15:0];
  assign nl_Product1_10_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5849:5845]));
  assign Product1_10_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6489:6485]));
  assign Product1_11_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_351_nl = (readslicef_20_16_4(Product1_10_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_351_nl = nl_Accum2_acc_351_nl[15:0];
  assign nl_Product1_12_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7129:7125]));
  assign Product1_12_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7769:7765]));
  assign Product1_13_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_350_nl = (readslicef_20_16_4(Product1_12_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_350_nl = nl_Accum2_acc_350_nl[15:0];
  assign nl_Accum2_acc_357_nl = Accum2_acc_351_nl + Accum2_acc_350_nl;
  assign Accum2_acc_357_nl = nl_Accum2_acc_357_nl[15:0];
  assign nl_Accum2_acc_1809_nl = (Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[89:85]);
  assign Accum2_acc_1809_nl = nl_Accum2_acc_1809_nl[9:0];
  assign nl_Product1_1_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[89:85]));
  assign Product1_1_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_356_nl = ({Accum2_acc_1809_nl , (Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_356_nl = nl_Accum2_acc_356_nl[15:0];
  assign nl_Accum2_acc_360_nl = Accum2_acc_357_nl + Accum2_acc_356_nl;
  assign Accum2_acc_360_nl = nl_Accum2_acc_360_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1 = Accum2_acc_361_nl
      + Accum2_acc_360_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[734:730]));
  assign Product1_2_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1374:1370]));
  assign Product1_3_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_368_nl = (readslicef_20_16_4(Product1_2_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_368_nl = nl_Accum2_acc_368_nl[15:0];
  assign nl_Product1_4_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2014:2010]));
  assign Product1_4_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2654:2650]));
  assign Product1_5_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_367_nl = (readslicef_20_16_4(Product1_4_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_367_nl = nl_Accum2_acc_367_nl[15:0];
  assign nl_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3294:3290]));
  assign Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3934:3930]));
  assign Product1_7_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_366_nl = (readslicef_20_16_4(Product1_6_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_366_nl = nl_Accum2_acc_366_nl[15:0];
  assign nl_Product1_8_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4574:4570]));
  assign Product1_8_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5214:5210]));
  assign Product1_9_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_365_nl = (readslicef_20_16_4(Product1_8_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_365_nl = nl_Accum2_acc_365_nl[15:0];
  assign nl_Accum2_acc_374_nl = Accum2_acc_368_nl + Accum2_acc_367_nl + Accum2_acc_366_nl
      + Accum2_acc_365_nl;
  assign Accum2_acc_374_nl = nl_Accum2_acc_374_nl[15:0];
  assign nl_Product1_10_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5854:5850]));
  assign Product1_10_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6494:6490]));
  assign Product1_11_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_364_nl = (readslicef_20_16_4(Product1_10_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_364_nl = nl_Accum2_acc_364_nl[15:0];
  assign nl_Product1_12_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7134:7130]));
  assign Product1_12_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7774:7770]));
  assign Product1_13_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_363_nl = (readslicef_20_16_4(Product1_12_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_363_nl = nl_Accum2_acc_363_nl[15:0];
  assign nl_Accum2_acc_370_nl = Accum2_acc_364_nl + Accum2_acc_363_nl;
  assign Accum2_acc_370_nl = nl_Accum2_acc_370_nl[15:0];
  assign nl_Accum2_acc_1810_nl = (Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[94:90]);
  assign Accum2_acc_1810_nl = nl_Accum2_acc_1810_nl[9:0];
  assign nl_Product1_1_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[94:90]));
  assign Product1_1_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_369_nl = ({Accum2_acc_1810_nl , (Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_369_nl = nl_Accum2_acc_369_nl[15:0];
  assign nl_Accum2_acc_373_nl = Accum2_acc_370_nl + Accum2_acc_369_nl;
  assign Accum2_acc_373_nl = nl_Accum2_acc_373_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1 = Accum2_acc_374_nl
      + Accum2_acc_373_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[739:735]));
  assign Product1_2_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1379:1375]));
  assign Product1_3_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_381_nl = (readslicef_20_16_4(Product1_2_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_381_nl = nl_Accum2_acc_381_nl[15:0];
  assign nl_Product1_4_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2019:2015]));
  assign Product1_4_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2659:2655]));
  assign Product1_5_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_380_nl = (readslicef_20_16_4(Product1_4_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_380_nl = nl_Accum2_acc_380_nl[15:0];
  assign nl_Product1_6_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3299:3295]));
  assign Product1_6_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3939:3935]));
  assign Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_379_nl = (readslicef_20_16_4(Product1_6_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_379_nl = nl_Accum2_acc_379_nl[15:0];
  assign nl_Product1_8_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4579:4575]));
  assign Product1_8_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5219:5215]));
  assign Product1_9_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_378_nl = (readslicef_20_16_4(Product1_8_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_378_nl = nl_Accum2_acc_378_nl[15:0];
  assign nl_Accum2_acc_387_nl = Accum2_acc_381_nl + Accum2_acc_380_nl + Accum2_acc_379_nl
      + Accum2_acc_378_nl;
  assign Accum2_acc_387_nl = nl_Accum2_acc_387_nl[15:0];
  assign nl_Product1_10_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5859:5855]));
  assign Product1_10_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6499:6495]));
  assign Product1_11_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_377_nl = (readslicef_20_16_4(Product1_10_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_377_nl = nl_Accum2_acc_377_nl[15:0];
  assign nl_Product1_12_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7139:7135]));
  assign Product1_12_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7779:7775]));
  assign Product1_13_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_376_nl = (readslicef_20_16_4(Product1_12_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_376_nl = nl_Accum2_acc_376_nl[15:0];
  assign nl_Accum2_acc_383_nl = Accum2_acc_377_nl + Accum2_acc_376_nl;
  assign Accum2_acc_383_nl = nl_Accum2_acc_383_nl[15:0];
  assign nl_Accum2_acc_1811_nl = (Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[99:95]);
  assign Accum2_acc_1811_nl = nl_Accum2_acc_1811_nl[9:0];
  assign nl_Product1_1_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[99:95]));
  assign Product1_1_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_382_nl = ({Accum2_acc_1811_nl , (Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_382_nl = nl_Accum2_acc_382_nl[15:0];
  assign nl_Accum2_acc_386_nl = Accum2_acc_383_nl + Accum2_acc_382_nl;
  assign Accum2_acc_386_nl = nl_Accum2_acc_386_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1 = Accum2_acc_387_nl
      + Accum2_acc_386_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[744:740]));
  assign Product1_2_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1384:1380]));
  assign Product1_3_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_394_nl = (readslicef_20_16_4(Product1_2_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_394_nl = nl_Accum2_acc_394_nl[15:0];
  assign nl_Product1_4_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2024:2020]));
  assign Product1_4_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2664:2660]));
  assign Product1_5_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_393_nl = (readslicef_20_16_4(Product1_4_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_393_nl = nl_Accum2_acc_393_nl[15:0];
  assign nl_Product1_6_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3304:3300]));
  assign Product1_6_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3944:3940]));
  assign Product1_7_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_392_nl = (readslicef_20_16_4(Product1_6_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_392_nl = nl_Accum2_acc_392_nl[15:0];
  assign nl_Product1_8_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4584:4580]));
  assign Product1_8_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5224:5220]));
  assign Product1_9_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_391_nl = (readslicef_20_16_4(Product1_8_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_391_nl = nl_Accum2_acc_391_nl[15:0];
  assign nl_Accum2_acc_400_nl = Accum2_acc_394_nl + Accum2_acc_393_nl + Accum2_acc_392_nl
      + Accum2_acc_391_nl;
  assign Accum2_acc_400_nl = nl_Accum2_acc_400_nl[15:0];
  assign nl_Product1_10_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5864:5860]));
  assign Product1_10_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6504:6500]));
  assign Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_390_nl = (readslicef_20_16_4(Product1_10_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_390_nl = nl_Accum2_acc_390_nl[15:0];
  assign nl_Product1_12_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7144:7140]));
  assign Product1_12_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7784:7780]));
  assign Product1_13_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_389_nl = (readslicef_20_16_4(Product1_12_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_389_nl = nl_Accum2_acc_389_nl[15:0];
  assign nl_Accum2_acc_396_nl = Accum2_acc_390_nl + Accum2_acc_389_nl;
  assign Accum2_acc_396_nl = nl_Accum2_acc_396_nl[15:0];
  assign nl_Accum2_acc_1812_nl = (Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[104:100]);
  assign Accum2_acc_1812_nl = nl_Accum2_acc_1812_nl[9:0];
  assign nl_Product1_1_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[104:100]));
  assign Product1_1_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_395_nl = ({Accum2_acc_1812_nl , (Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_395_nl = nl_Accum2_acc_395_nl[15:0];
  assign nl_Accum2_acc_399_nl = Accum2_acc_396_nl + Accum2_acc_395_nl;
  assign Accum2_acc_399_nl = nl_Accum2_acc_399_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1 = Accum2_acc_400_nl
      + Accum2_acc_399_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[749:745]));
  assign Product1_2_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1389:1385]));
  assign Product1_3_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_407_nl = (readslicef_20_16_4(Product1_2_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_407_nl = nl_Accum2_acc_407_nl[15:0];
  assign nl_Product1_4_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2029:2025]));
  assign Product1_4_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2669:2665]));
  assign Product1_5_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_406_nl = (readslicef_20_16_4(Product1_4_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_406_nl = nl_Accum2_acc_406_nl[15:0];
  assign nl_Product1_6_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3309:3305]));
  assign Product1_6_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3949:3945]));
  assign Product1_7_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_405_nl = (readslicef_20_16_4(Product1_6_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_405_nl = nl_Accum2_acc_405_nl[15:0];
  assign nl_Product1_8_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4589:4585]));
  assign Product1_8_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5229:5225]));
  assign Product1_9_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_404_nl = (readslicef_20_16_4(Product1_8_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_404_nl = nl_Accum2_acc_404_nl[15:0];
  assign nl_Accum2_acc_413_nl = Accum2_acc_407_nl + Accum2_acc_406_nl + Accum2_acc_405_nl
      + Accum2_acc_404_nl;
  assign Accum2_acc_413_nl = nl_Accum2_acc_413_nl[15:0];
  assign nl_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5869:5865]));
  assign Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6509:6505]));
  assign Product1_11_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_403_nl = (readslicef_20_16_4(Product1_10_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_403_nl = nl_Accum2_acc_403_nl[15:0];
  assign nl_Product1_12_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7149:7145]));
  assign Product1_12_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7789:7785]));
  assign Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_402_nl = (readslicef_20_16_4(Product1_12_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_402_nl = nl_Accum2_acc_402_nl[15:0];
  assign nl_Accum2_acc_409_nl = Accum2_acc_403_nl + Accum2_acc_402_nl;
  assign Accum2_acc_409_nl = nl_Accum2_acc_409_nl[15:0];
  assign nl_Accum2_acc_1813_nl = (Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[109:105]);
  assign Accum2_acc_1813_nl = nl_Accum2_acc_1813_nl[9:0];
  assign nl_Product1_1_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[109:105]));
  assign Product1_1_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_408_nl = ({Accum2_acc_1813_nl , (Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_408_nl = nl_Accum2_acc_408_nl[15:0];
  assign nl_Accum2_acc_412_nl = Accum2_acc_409_nl + Accum2_acc_408_nl;
  assign Accum2_acc_412_nl = nl_Accum2_acc_412_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1 = Accum2_acc_413_nl
      + Accum2_acc_412_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[754:750]));
  assign Product1_2_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1394:1390]));
  assign Product1_3_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_420_nl = (readslicef_20_16_4(Product1_2_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_420_nl = nl_Accum2_acc_420_nl[15:0];
  assign nl_Product1_4_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2034:2030]));
  assign Product1_4_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2674:2670]));
  assign Product1_5_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_419_nl = (readslicef_20_16_4(Product1_4_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_419_nl = nl_Accum2_acc_419_nl[15:0];
  assign nl_Product1_6_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3314:3310]));
  assign Product1_6_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3954:3950]));
  assign Product1_7_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_418_nl = (readslicef_20_16_4(Product1_6_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_418_nl = nl_Accum2_acc_418_nl[15:0];
  assign nl_Product1_8_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4594:4590]));
  assign Product1_8_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5234:5230]));
  assign Product1_9_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_417_nl = (readslicef_20_16_4(Product1_8_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_417_nl = nl_Accum2_acc_417_nl[15:0];
  assign nl_Accum2_acc_426_nl = Accum2_acc_420_nl + Accum2_acc_419_nl + Accum2_acc_418_nl
      + Accum2_acc_417_nl;
  assign Accum2_acc_426_nl = nl_Accum2_acc_426_nl[15:0];
  assign nl_Product1_10_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5874:5870]));
  assign Product1_10_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6514:6510]));
  assign Product1_11_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_416_nl = (readslicef_20_16_4(Product1_10_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_416_nl = nl_Accum2_acc_416_nl[15:0];
  assign nl_Product1_12_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7154:7150]));
  assign Product1_12_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7794:7790]));
  assign Product1_13_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_415_nl = (readslicef_20_16_4(Product1_12_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_415_nl = nl_Accum2_acc_415_nl[15:0];
  assign nl_Accum2_acc_422_nl = Accum2_acc_416_nl + Accum2_acc_415_nl;
  assign Accum2_acc_422_nl = nl_Accum2_acc_422_nl[15:0];
  assign nl_Accum2_acc_1814_nl = (Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[114:110]);
  assign Accum2_acc_1814_nl = nl_Accum2_acc_1814_nl[9:0];
  assign nl_Product1_1_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[114:110]));
  assign Product1_1_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_421_nl = ({Accum2_acc_1814_nl , (Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_421_nl = nl_Accum2_acc_421_nl[15:0];
  assign nl_Accum2_acc_425_nl = Accum2_acc_422_nl + Accum2_acc_421_nl;
  assign Accum2_acc_425_nl = nl_Accum2_acc_425_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1 = Accum2_acc_426_nl
      + Accum2_acc_425_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[759:755]));
  assign Product1_2_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1399:1395]));
  assign Product1_3_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_433_nl = (readslicef_20_16_4(Product1_2_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_433_nl = nl_Accum2_acc_433_nl[15:0];
  assign nl_Product1_4_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2039:2035]));
  assign Product1_4_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2679:2675]));
  assign Product1_5_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_432_nl = (readslicef_20_16_4(Product1_4_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_432_nl = nl_Accum2_acc_432_nl[15:0];
  assign nl_Product1_6_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3319:3315]));
  assign Product1_6_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3959:3955]));
  assign Product1_7_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_431_nl = (readslicef_20_16_4(Product1_6_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_431_nl = nl_Accum2_acc_431_nl[15:0];
  assign nl_Product1_8_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4599:4595]));
  assign Product1_8_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5239:5235]));
  assign Product1_9_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_430_nl = (readslicef_20_16_4(Product1_8_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_430_nl = nl_Accum2_acc_430_nl[15:0];
  assign nl_Accum2_acc_439_nl = Accum2_acc_433_nl + Accum2_acc_432_nl + Accum2_acc_431_nl
      + Accum2_acc_430_nl;
  assign Accum2_acc_439_nl = nl_Accum2_acc_439_nl[15:0];
  assign nl_Product1_10_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5879:5875]));
  assign Product1_10_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6519:6515]));
  assign Product1_11_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_429_nl = (readslicef_20_16_4(Product1_10_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_429_nl = nl_Accum2_acc_429_nl[15:0];
  assign nl_Product1_12_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7159:7155]));
  assign Product1_12_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7799:7795]));
  assign Product1_13_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_428_nl = (readslicef_20_16_4(Product1_12_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_428_nl = nl_Accum2_acc_428_nl[15:0];
  assign nl_Accum2_acc_435_nl = Accum2_acc_429_nl + Accum2_acc_428_nl;
  assign Accum2_acc_435_nl = nl_Accum2_acc_435_nl[15:0];
  assign nl_Accum2_acc_1815_nl = (Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[119:115]);
  assign Accum2_acc_1815_nl = nl_Accum2_acc_1815_nl[9:0];
  assign nl_Product1_1_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[119:115]));
  assign Product1_1_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_434_nl = ({Accum2_acc_1815_nl , (Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_434_nl = nl_Accum2_acc_434_nl[15:0];
  assign nl_Accum2_acc_438_nl = Accum2_acc_435_nl + Accum2_acc_434_nl;
  assign Accum2_acc_438_nl = nl_Accum2_acc_438_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1 = Accum2_acc_439_nl
      + Accum2_acc_438_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[764:760]));
  assign Product1_2_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1404:1400]));
  assign Product1_3_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_446_nl = (readslicef_20_16_4(Product1_2_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_446_nl = nl_Accum2_acc_446_nl[15:0];
  assign nl_Product1_4_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2044:2040]));
  assign Product1_4_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2684:2680]));
  assign Product1_5_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_445_nl = (readslicef_20_16_4(Product1_4_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_445_nl = nl_Accum2_acc_445_nl[15:0];
  assign nl_Product1_6_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3324:3320]));
  assign Product1_6_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3964:3960]));
  assign Product1_7_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_444_nl = (readslicef_20_16_4(Product1_6_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_444_nl = nl_Accum2_acc_444_nl[15:0];
  assign nl_Product1_8_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4604:4600]));
  assign Product1_8_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5244:5240]));
  assign Product1_9_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_443_nl = (readslicef_20_16_4(Product1_8_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_443_nl = nl_Accum2_acc_443_nl[15:0];
  assign nl_Accum2_acc_452_nl = Accum2_acc_446_nl + Accum2_acc_445_nl + Accum2_acc_444_nl
      + Accum2_acc_443_nl;
  assign Accum2_acc_452_nl = nl_Accum2_acc_452_nl[15:0];
  assign nl_Product1_10_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5884:5880]));
  assign Product1_10_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6524:6520]));
  assign Product1_11_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_442_nl = (readslicef_20_16_4(Product1_10_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_442_nl = nl_Accum2_acc_442_nl[15:0];
  assign nl_Product1_12_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7164:7160]));
  assign Product1_12_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7804:7800]));
  assign Product1_13_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_441_nl = (readslicef_20_16_4(Product1_12_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_441_nl = nl_Accum2_acc_441_nl[15:0];
  assign nl_Accum2_acc_448_nl = Accum2_acc_442_nl + Accum2_acc_441_nl;
  assign Accum2_acc_448_nl = nl_Accum2_acc_448_nl[15:0];
  assign nl_Accum2_acc_1816_nl = (Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[124:120]);
  assign Accum2_acc_1816_nl = nl_Accum2_acc_1816_nl[9:0];
  assign nl_Product1_1_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[124:120]));
  assign Product1_1_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_447_nl = ({Accum2_acc_1816_nl , (Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_447_nl = nl_Accum2_acc_447_nl[15:0];
  assign nl_Accum2_acc_451_nl = Accum2_acc_448_nl + Accum2_acc_447_nl;
  assign Accum2_acc_451_nl = nl_Accum2_acc_451_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1 = Accum2_acc_452_nl
      + Accum2_acc_451_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[769:765]));
  assign Product1_2_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1409:1405]));
  assign Product1_3_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_459_nl = (readslicef_20_16_4(Product1_2_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_459_nl = nl_Accum2_acc_459_nl[15:0];
  assign nl_Product1_4_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2049:2045]));
  assign Product1_4_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2689:2685]));
  assign Product1_5_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_458_nl = (readslicef_20_16_4(Product1_4_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_458_nl = nl_Accum2_acc_458_nl[15:0];
  assign nl_Product1_6_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3329:3325]));
  assign Product1_6_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3969:3965]));
  assign Product1_7_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_457_nl = (readslicef_20_16_4(Product1_6_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_457_nl = nl_Accum2_acc_457_nl[15:0];
  assign nl_Product1_8_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4609:4605]));
  assign Product1_8_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5249:5245]));
  assign Product1_9_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_456_nl = (readslicef_20_16_4(Product1_8_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_456_nl = nl_Accum2_acc_456_nl[15:0];
  assign nl_Accum2_acc_465_nl = Accum2_acc_459_nl + Accum2_acc_458_nl + Accum2_acc_457_nl
      + Accum2_acc_456_nl;
  assign Accum2_acc_465_nl = nl_Accum2_acc_465_nl[15:0];
  assign nl_Product1_10_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5889:5885]));
  assign Product1_10_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6529:6525]));
  assign Product1_11_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_455_nl = (readslicef_20_16_4(Product1_10_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_455_nl = nl_Accum2_acc_455_nl[15:0];
  assign nl_Product1_12_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7169:7165]));
  assign Product1_12_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7809:7805]));
  assign Product1_13_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_454_nl = (readslicef_20_16_4(Product1_12_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_454_nl = nl_Accum2_acc_454_nl[15:0];
  assign nl_Accum2_acc_461_nl = Accum2_acc_455_nl + Accum2_acc_454_nl;
  assign Accum2_acc_461_nl = nl_Accum2_acc_461_nl[15:0];
  assign nl_Accum2_acc_1817_nl = (Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[129:125]);
  assign Accum2_acc_1817_nl = nl_Accum2_acc_1817_nl[9:0];
  assign nl_Product1_1_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[129:125]));
  assign Product1_1_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_460_nl = ({Accum2_acc_1817_nl , (Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_460_nl = nl_Accum2_acc_460_nl[15:0];
  assign nl_Accum2_acc_464_nl = Accum2_acc_461_nl + Accum2_acc_460_nl;
  assign Accum2_acc_464_nl = nl_Accum2_acc_464_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1 = Accum2_acc_465_nl
      + Accum2_acc_464_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[774:770]));
  assign Product1_2_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1414:1410]));
  assign Product1_3_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_472_nl = (readslicef_20_16_4(Product1_2_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_472_nl = nl_Accum2_acc_472_nl[15:0];
  assign nl_Product1_4_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2054:2050]));
  assign Product1_4_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2694:2690]));
  assign Product1_5_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_471_nl = (readslicef_20_16_4(Product1_4_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_471_nl = nl_Accum2_acc_471_nl[15:0];
  assign nl_Product1_6_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3334:3330]));
  assign Product1_6_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3974:3970]));
  assign Product1_7_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_470_nl = (readslicef_20_16_4(Product1_6_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_470_nl = nl_Accum2_acc_470_nl[15:0];
  assign nl_Product1_8_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4614:4610]));
  assign Product1_8_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5254:5250]));
  assign Product1_9_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_469_nl = (readslicef_20_16_4(Product1_8_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_469_nl = nl_Accum2_acc_469_nl[15:0];
  assign nl_Accum2_acc_478_nl = Accum2_acc_472_nl + Accum2_acc_471_nl + Accum2_acc_470_nl
      + Accum2_acc_469_nl;
  assign Accum2_acc_478_nl = nl_Accum2_acc_478_nl[15:0];
  assign nl_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5894:5890]));
  assign Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6534:6530]));
  assign Product1_11_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_468_nl = (readslicef_20_16_4(Product1_10_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_468_nl = nl_Accum2_acc_468_nl[15:0];
  assign nl_Product1_12_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7174:7170]));
  assign Product1_12_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7814:7810]));
  assign Product1_13_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_467_nl = (readslicef_20_16_4(Product1_12_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_467_nl = nl_Accum2_acc_467_nl[15:0];
  assign nl_Accum2_acc_474_nl = Accum2_acc_468_nl + Accum2_acc_467_nl;
  assign Accum2_acc_474_nl = nl_Accum2_acc_474_nl[15:0];
  assign nl_Accum2_acc_1818_nl = (Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[134:130]);
  assign Accum2_acc_1818_nl = nl_Accum2_acc_1818_nl[9:0];
  assign nl_Product1_1_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[134:130]));
  assign Product1_1_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_473_nl = ({Accum2_acc_1818_nl , (Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_473_nl = nl_Accum2_acc_473_nl[15:0];
  assign nl_Accum2_acc_477_nl = Accum2_acc_474_nl + Accum2_acc_473_nl;
  assign Accum2_acc_477_nl = nl_Accum2_acc_477_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1 = Accum2_acc_478_nl
      + Accum2_acc_477_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[779:775]));
  assign Product1_2_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1419:1415]));
  assign Product1_3_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_485_nl = (readslicef_20_16_4(Product1_2_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_485_nl = nl_Accum2_acc_485_nl[15:0];
  assign nl_Product1_4_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2059:2055]));
  assign Product1_4_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2699:2695]));
  assign Product1_5_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_484_nl = (readslicef_20_16_4(Product1_4_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_484_nl = nl_Accum2_acc_484_nl[15:0];
  assign nl_Product1_6_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3339:3335]));
  assign Product1_6_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3979:3975]));
  assign Product1_7_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_483_nl = (readslicef_20_16_4(Product1_6_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_483_nl = nl_Accum2_acc_483_nl[15:0];
  assign nl_Product1_8_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4619:4615]));
  assign Product1_8_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5259:5255]));
  assign Product1_9_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_482_nl = (readslicef_20_16_4(Product1_8_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_482_nl = nl_Accum2_acc_482_nl[15:0];
  assign nl_Accum2_acc_491_nl = Accum2_acc_485_nl + Accum2_acc_484_nl + Accum2_acc_483_nl
      + Accum2_acc_482_nl;
  assign Accum2_acc_491_nl = nl_Accum2_acc_491_nl[15:0];
  assign nl_Product1_10_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5899:5895]));
  assign Product1_10_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6539:6535]));
  assign Product1_11_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_481_nl = (readslicef_20_16_4(Product1_10_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_481_nl = nl_Accum2_acc_481_nl[15:0];
  assign nl_Product1_12_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7179:7175]));
  assign Product1_12_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7819:7815]));
  assign Product1_13_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_480_nl = (readslicef_20_16_4(Product1_12_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_480_nl = nl_Accum2_acc_480_nl[15:0];
  assign nl_Accum2_acc_487_nl = Accum2_acc_481_nl + Accum2_acc_480_nl;
  assign Accum2_acc_487_nl = nl_Accum2_acc_487_nl[15:0];
  assign nl_Accum2_acc_1819_nl = (Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[139:135]);
  assign Accum2_acc_1819_nl = nl_Accum2_acc_1819_nl[9:0];
  assign nl_Product1_1_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[139:135]));
  assign Product1_1_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_486_nl = ({Accum2_acc_1819_nl , (Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_486_nl = nl_Accum2_acc_486_nl[15:0];
  assign nl_Accum2_acc_490_nl = Accum2_acc_487_nl + Accum2_acc_486_nl;
  assign Accum2_acc_490_nl = nl_Accum2_acc_490_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1 = Accum2_acc_491_nl
      + Accum2_acc_490_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[784:780]));
  assign Product1_2_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1424:1420]));
  assign Product1_3_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_498_nl = (readslicef_20_16_4(Product1_2_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_498_nl = nl_Accum2_acc_498_nl[15:0];
  assign nl_Product1_4_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2064:2060]));
  assign Product1_4_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2704:2700]));
  assign Product1_5_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_497_nl = (readslicef_20_16_4(Product1_4_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_497_nl = nl_Accum2_acc_497_nl[15:0];
  assign nl_Product1_6_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3344:3340]));
  assign Product1_6_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3984:3980]));
  assign Product1_7_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_496_nl = (readslicef_20_16_4(Product1_6_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_496_nl = nl_Accum2_acc_496_nl[15:0];
  assign nl_Product1_8_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4624:4620]));
  assign Product1_8_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5264:5260]));
  assign Product1_9_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_495_nl = (readslicef_20_16_4(Product1_8_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_495_nl = nl_Accum2_acc_495_nl[15:0];
  assign nl_Accum2_acc_504_nl = Accum2_acc_498_nl + Accum2_acc_497_nl + Accum2_acc_496_nl
      + Accum2_acc_495_nl;
  assign Accum2_acc_504_nl = nl_Accum2_acc_504_nl[15:0];
  assign nl_Product1_10_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5904:5900]));
  assign Product1_10_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6544:6540]));
  assign Product1_11_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_494_nl = (readslicef_20_16_4(Product1_10_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_494_nl = nl_Accum2_acc_494_nl[15:0];
  assign nl_Product1_12_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7184:7180]));
  assign Product1_12_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7824:7820]));
  assign Product1_13_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_493_nl = (readslicef_20_16_4(Product1_12_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_493_nl = nl_Accum2_acc_493_nl[15:0];
  assign nl_Accum2_acc_500_nl = Accum2_acc_494_nl + Accum2_acc_493_nl;
  assign Accum2_acc_500_nl = nl_Accum2_acc_500_nl[15:0];
  assign nl_Accum2_acc_1820_nl = (Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[144:140]);
  assign Accum2_acc_1820_nl = nl_Accum2_acc_1820_nl[9:0];
  assign nl_Product1_1_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[144:140]));
  assign Product1_1_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_499_nl = ({Accum2_acc_1820_nl , (Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_499_nl = nl_Accum2_acc_499_nl[15:0];
  assign nl_Accum2_acc_503_nl = Accum2_acc_500_nl + Accum2_acc_499_nl;
  assign Accum2_acc_503_nl = nl_Accum2_acc_503_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1 = Accum2_acc_504_nl
      + Accum2_acc_503_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[789:785]));
  assign Product1_2_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1429:1425]));
  assign Product1_3_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_511_nl = (readslicef_20_16_4(Product1_2_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_511_nl = nl_Accum2_acc_511_nl[15:0];
  assign nl_Product1_4_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2069:2065]));
  assign Product1_4_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2709:2705]));
  assign Product1_5_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_510_nl = (readslicef_20_16_4(Product1_4_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_510_nl = nl_Accum2_acc_510_nl[15:0];
  assign nl_Product1_6_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3349:3345]));
  assign Product1_6_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3989:3985]));
  assign Product1_7_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_509_nl = (readslicef_20_16_4(Product1_6_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_509_nl = nl_Accum2_acc_509_nl[15:0];
  assign nl_Product1_8_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4629:4625]));
  assign Product1_8_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5269:5265]));
  assign Product1_9_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_508_nl = (readslicef_20_16_4(Product1_8_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_508_nl = nl_Accum2_acc_508_nl[15:0];
  assign nl_Accum2_acc_517_nl = Accum2_acc_511_nl + Accum2_acc_510_nl + Accum2_acc_509_nl
      + Accum2_acc_508_nl;
  assign Accum2_acc_517_nl = nl_Accum2_acc_517_nl[15:0];
  assign nl_Product1_10_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5909:5905]));
  assign Product1_10_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6549:6545]));
  assign Product1_11_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_507_nl = (readslicef_20_16_4(Product1_10_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_507_nl = nl_Accum2_acc_507_nl[15:0];
  assign nl_Product1_12_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7189:7185]));
  assign Product1_12_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7829:7825]));
  assign Product1_13_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_506_nl = (readslicef_20_16_4(Product1_12_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_506_nl = nl_Accum2_acc_506_nl[15:0];
  assign nl_Accum2_acc_513_nl = Accum2_acc_507_nl + Accum2_acc_506_nl;
  assign Accum2_acc_513_nl = nl_Accum2_acc_513_nl[15:0];
  assign nl_Accum2_acc_1821_nl = (Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[149:145]);
  assign Accum2_acc_1821_nl = nl_Accum2_acc_1821_nl[9:0];
  assign nl_Product1_1_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[149:145]));
  assign Product1_1_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_512_nl = ({Accum2_acc_1821_nl , (Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_512_nl = nl_Accum2_acc_512_nl[15:0];
  assign nl_Accum2_acc_516_nl = Accum2_acc_513_nl + Accum2_acc_512_nl;
  assign Accum2_acc_516_nl = nl_Accum2_acc_516_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1 = Accum2_acc_517_nl
      + Accum2_acc_516_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[794:790]));
  assign Product1_2_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1434:1430]));
  assign Product1_3_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_524_nl = (readslicef_20_16_4(Product1_2_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_524_nl = nl_Accum2_acc_524_nl[15:0];
  assign nl_Product1_4_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2074:2070]));
  assign Product1_4_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2714:2710]));
  assign Product1_5_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_523_nl = (readslicef_20_16_4(Product1_4_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_523_nl = nl_Accum2_acc_523_nl[15:0];
  assign nl_Product1_6_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3354:3350]));
  assign Product1_6_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3994:3990]));
  assign Product1_7_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_522_nl = (readslicef_20_16_4(Product1_6_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_522_nl = nl_Accum2_acc_522_nl[15:0];
  assign nl_Product1_8_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4634:4630]));
  assign Product1_8_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5274:5270]));
  assign Product1_9_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_521_nl = (readslicef_20_16_4(Product1_8_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_521_nl = nl_Accum2_acc_521_nl[15:0];
  assign nl_Accum2_acc_530_nl = Accum2_acc_524_nl + Accum2_acc_523_nl + Accum2_acc_522_nl
      + Accum2_acc_521_nl;
  assign Accum2_acc_530_nl = nl_Accum2_acc_530_nl[15:0];
  assign nl_Product1_10_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5914:5910]));
  assign Product1_10_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6554:6550]));
  assign Product1_11_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_520_nl = (readslicef_20_16_4(Product1_10_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_520_nl = nl_Accum2_acc_520_nl[15:0];
  assign nl_Product1_12_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7194:7190]));
  assign Product1_12_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7834:7830]));
  assign Product1_13_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_519_nl = (readslicef_20_16_4(Product1_12_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_519_nl = nl_Accum2_acc_519_nl[15:0];
  assign nl_Accum2_acc_526_nl = Accum2_acc_520_nl + Accum2_acc_519_nl;
  assign Accum2_acc_526_nl = nl_Accum2_acc_526_nl[15:0];
  assign nl_Accum2_acc_1822_nl = (Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[154:150]);
  assign Accum2_acc_1822_nl = nl_Accum2_acc_1822_nl[9:0];
  assign nl_Product1_1_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[154:150]));
  assign Product1_1_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_525_nl = ({Accum2_acc_1822_nl , (Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_525_nl = nl_Accum2_acc_525_nl[15:0];
  assign nl_Accum2_acc_529_nl = Accum2_acc_526_nl + Accum2_acc_525_nl;
  assign Accum2_acc_529_nl = nl_Accum2_acc_529_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1 = Accum2_acc_530_nl
      + Accum2_acc_529_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[799:795]));
  assign Product1_2_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1439:1435]));
  assign Product1_3_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_537_nl = (readslicef_20_16_4(Product1_2_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_537_nl = nl_Accum2_acc_537_nl[15:0];
  assign nl_Product1_4_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2079:2075]));
  assign Product1_4_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2719:2715]));
  assign Product1_5_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_536_nl = (readslicef_20_16_4(Product1_4_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_536_nl = nl_Accum2_acc_536_nl[15:0];
  assign nl_Product1_6_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3359:3355]));
  assign Product1_6_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[3999:3995]));
  assign Product1_7_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_535_nl = (readslicef_20_16_4(Product1_6_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_535_nl = nl_Accum2_acc_535_nl[15:0];
  assign nl_Product1_8_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4639:4635]));
  assign Product1_8_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5279:5275]));
  assign Product1_9_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_534_nl = (readslicef_20_16_4(Product1_8_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_534_nl = nl_Accum2_acc_534_nl[15:0];
  assign nl_Accum2_acc_543_nl = Accum2_acc_537_nl + Accum2_acc_536_nl + Accum2_acc_535_nl
      + Accum2_acc_534_nl;
  assign Accum2_acc_543_nl = nl_Accum2_acc_543_nl[15:0];
  assign nl_Product1_10_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5919:5915]));
  assign Product1_10_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6559:6555]));
  assign Product1_11_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_533_nl = (readslicef_20_16_4(Product1_10_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_533_nl = nl_Accum2_acc_533_nl[15:0];
  assign nl_Product1_12_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7199:7195]));
  assign Product1_12_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7839:7835]));
  assign Product1_13_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_532_nl = (readslicef_20_16_4(Product1_12_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_532_nl = nl_Accum2_acc_532_nl[15:0];
  assign nl_Accum2_acc_539_nl = Accum2_acc_533_nl + Accum2_acc_532_nl;
  assign Accum2_acc_539_nl = nl_Accum2_acc_539_nl[15:0];
  assign nl_Accum2_acc_1823_nl = (Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[159:155]);
  assign Accum2_acc_1823_nl = nl_Accum2_acc_1823_nl[9:0];
  assign nl_Product1_1_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[159:155]));
  assign Product1_1_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_538_nl = ({Accum2_acc_1823_nl , (Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_538_nl = nl_Accum2_acc_538_nl[15:0];
  assign nl_Accum2_acc_542_nl = Accum2_acc_539_nl + Accum2_acc_538_nl;
  assign Accum2_acc_542_nl = nl_Accum2_acc_542_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1 = Accum2_acc_543_nl
      + Accum2_acc_542_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[804:800]));
  assign Product1_2_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1444:1440]));
  assign Product1_3_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_550_nl = (readslicef_20_16_4(Product1_2_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_550_nl = nl_Accum2_acc_550_nl[15:0];
  assign nl_Product1_4_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2084:2080]));
  assign Product1_4_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2724:2720]));
  assign Product1_5_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_549_nl = (readslicef_20_16_4(Product1_4_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_549_nl = nl_Accum2_acc_549_nl[15:0];
  assign nl_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3364:3360]));
  assign Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4004:4000]));
  assign Product1_7_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_548_nl = (readslicef_20_16_4(Product1_6_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_548_nl = nl_Accum2_acc_548_nl[15:0];
  assign nl_Product1_8_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4644:4640]));
  assign Product1_8_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5284:5280]));
  assign Product1_9_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_547_nl = (readslicef_20_16_4(Product1_8_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_547_nl = nl_Accum2_acc_547_nl[15:0];
  assign nl_Accum2_acc_556_nl = Accum2_acc_550_nl + Accum2_acc_549_nl + Accum2_acc_548_nl
      + Accum2_acc_547_nl;
  assign Accum2_acc_556_nl = nl_Accum2_acc_556_nl[15:0];
  assign nl_Product1_10_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5924:5920]));
  assign Product1_10_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6564:6560]));
  assign Product1_11_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_546_nl = (readslicef_20_16_4(Product1_10_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_546_nl = nl_Accum2_acc_546_nl[15:0];
  assign nl_Product1_12_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7204:7200]));
  assign Product1_12_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7844:7840]));
  assign Product1_13_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_545_nl = (readslicef_20_16_4(Product1_12_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_545_nl = nl_Accum2_acc_545_nl[15:0];
  assign nl_Accum2_acc_552_nl = Accum2_acc_546_nl + Accum2_acc_545_nl;
  assign Accum2_acc_552_nl = nl_Accum2_acc_552_nl[15:0];
  assign nl_Accum2_acc_1824_nl = (Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[164:160]);
  assign Accum2_acc_1824_nl = nl_Accum2_acc_1824_nl[9:0];
  assign nl_Product1_1_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[164:160]));
  assign Product1_1_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_551_nl = ({Accum2_acc_1824_nl , (Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_551_nl = nl_Accum2_acc_551_nl[15:0];
  assign nl_Accum2_acc_555_nl = Accum2_acc_552_nl + Accum2_acc_551_nl;
  assign Accum2_acc_555_nl = nl_Accum2_acc_555_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1 = Accum2_acc_556_nl
      + Accum2_acc_555_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[809:805]));
  assign Product1_2_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1449:1445]));
  assign Product1_3_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_563_nl = (readslicef_20_16_4(Product1_2_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_563_nl = nl_Accum2_acc_563_nl[15:0];
  assign nl_Product1_4_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2089:2085]));
  assign Product1_4_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2729:2725]));
  assign Product1_5_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_562_nl = (readslicef_20_16_4(Product1_4_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_562_nl = nl_Accum2_acc_562_nl[15:0];
  assign nl_Product1_6_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3369:3365]));
  assign Product1_6_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4009:4005]));
  assign Product1_7_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_561_nl = (readslicef_20_16_4(Product1_6_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_561_nl = nl_Accum2_acc_561_nl[15:0];
  assign nl_Product1_8_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4649:4645]));
  assign Product1_8_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5289:5285]));
  assign Product1_9_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_560_nl = (readslicef_20_16_4(Product1_8_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_560_nl = nl_Accum2_acc_560_nl[15:0];
  assign nl_Accum2_acc_569_nl = Accum2_acc_563_nl + Accum2_acc_562_nl + Accum2_acc_561_nl
      + Accum2_acc_560_nl;
  assign Accum2_acc_569_nl = nl_Accum2_acc_569_nl[15:0];
  assign nl_Product1_10_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5929:5925]));
  assign Product1_10_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6569:6565]));
  assign Product1_11_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_559_nl = (readslicef_20_16_4(Product1_10_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_559_nl = nl_Accum2_acc_559_nl[15:0];
  assign nl_Product1_12_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7209:7205]));
  assign Product1_12_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7849:7845]));
  assign Product1_13_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_558_nl = (readslicef_20_16_4(Product1_12_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_558_nl = nl_Accum2_acc_558_nl[15:0];
  assign nl_Accum2_acc_565_nl = Accum2_acc_559_nl + Accum2_acc_558_nl;
  assign Accum2_acc_565_nl = nl_Accum2_acc_565_nl[15:0];
  assign nl_Accum2_acc_1825_nl = (Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[169:165]);
  assign Accum2_acc_1825_nl = nl_Accum2_acc_1825_nl[9:0];
  assign nl_Product1_1_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[169:165]));
  assign Product1_1_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_564_nl = ({Accum2_acc_1825_nl , (Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_564_nl = nl_Accum2_acc_564_nl[15:0];
  assign nl_Accum2_acc_568_nl = Accum2_acc_565_nl + Accum2_acc_564_nl;
  assign Accum2_acc_568_nl = nl_Accum2_acc_568_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1 = Accum2_acc_569_nl
      + Accum2_acc_568_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[814:810]));
  assign Product1_2_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1454:1450]));
  assign Product1_3_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_576_nl = (readslicef_20_16_4(Product1_2_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_576_nl = nl_Accum2_acc_576_nl[15:0];
  assign nl_Product1_4_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2094:2090]));
  assign Product1_4_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2734:2730]));
  assign Product1_5_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_575_nl = (readslicef_20_16_4(Product1_4_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_575_nl = nl_Accum2_acc_575_nl[15:0];
  assign nl_Product1_6_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3374:3370]));
  assign Product1_6_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4014:4010]));
  assign Product1_7_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_574_nl = (readslicef_20_16_4(Product1_6_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_574_nl = nl_Accum2_acc_574_nl[15:0];
  assign nl_Product1_8_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4654:4650]));
  assign Product1_8_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5294:5290]));
  assign Product1_9_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_573_nl = (readslicef_20_16_4(Product1_8_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_573_nl = nl_Accum2_acc_573_nl[15:0];
  assign nl_Accum2_acc_582_nl = Accum2_acc_576_nl + Accum2_acc_575_nl + Accum2_acc_574_nl
      + Accum2_acc_573_nl;
  assign Accum2_acc_582_nl = nl_Accum2_acc_582_nl[15:0];
  assign nl_Product1_10_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5934:5930]));
  assign Product1_10_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6574:6570]));
  assign Product1_11_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_572_nl = (readslicef_20_16_4(Product1_10_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_572_nl = nl_Accum2_acc_572_nl[15:0];
  assign nl_Product1_12_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7214:7210]));
  assign Product1_12_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7854:7850]));
  assign Product1_13_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_571_nl = (readslicef_20_16_4(Product1_12_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_571_nl = nl_Accum2_acc_571_nl[15:0];
  assign nl_Accum2_acc_578_nl = Accum2_acc_572_nl + Accum2_acc_571_nl;
  assign Accum2_acc_578_nl = nl_Accum2_acc_578_nl[15:0];
  assign nl_Accum2_acc_1826_nl = (Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[174:170]);
  assign Accum2_acc_1826_nl = nl_Accum2_acc_1826_nl[9:0];
  assign nl_Product1_1_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[174:170]));
  assign Product1_1_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_577_nl = ({Accum2_acc_1826_nl , (Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_577_nl = nl_Accum2_acc_577_nl[15:0];
  assign nl_Accum2_acc_581_nl = Accum2_acc_578_nl + Accum2_acc_577_nl;
  assign Accum2_acc_581_nl = nl_Accum2_acc_581_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1 = Accum2_acc_582_nl
      + Accum2_acc_581_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[819:815]));
  assign Product1_2_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1459:1455]));
  assign Product1_3_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_589_nl = (readslicef_20_16_4(Product1_2_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_589_nl = nl_Accum2_acc_589_nl[15:0];
  assign nl_Product1_4_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2099:2095]));
  assign Product1_4_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2739:2735]));
  assign Product1_5_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_588_nl = (readslicef_20_16_4(Product1_4_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_588_nl = nl_Accum2_acc_588_nl[15:0];
  assign nl_Product1_6_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3379:3375]));
  assign Product1_6_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4019:4015]));
  assign Product1_7_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_587_nl = (readslicef_20_16_4(Product1_6_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_587_nl = nl_Accum2_acc_587_nl[15:0];
  assign nl_Product1_8_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4659:4655]));
  assign Product1_8_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5299:5295]));
  assign Product1_9_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_586_nl = (readslicef_20_16_4(Product1_8_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_586_nl = nl_Accum2_acc_586_nl[15:0];
  assign nl_Accum2_acc_595_nl = Accum2_acc_589_nl + Accum2_acc_588_nl + Accum2_acc_587_nl
      + Accum2_acc_586_nl;
  assign Accum2_acc_595_nl = nl_Accum2_acc_595_nl[15:0];
  assign nl_Product1_10_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5939:5935]));
  assign Product1_10_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6579:6575]));
  assign Product1_11_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_585_nl = (readslicef_20_16_4(Product1_10_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_585_nl = nl_Accum2_acc_585_nl[15:0];
  assign nl_Product1_12_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7219:7215]));
  assign Product1_12_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7859:7855]));
  assign Product1_13_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_584_nl = (readslicef_20_16_4(Product1_12_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_584_nl = nl_Accum2_acc_584_nl[15:0];
  assign nl_Accum2_acc_591_nl = Accum2_acc_585_nl + Accum2_acc_584_nl;
  assign Accum2_acc_591_nl = nl_Accum2_acc_591_nl[15:0];
  assign nl_Accum2_acc_1827_nl = (Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[179:175]);
  assign Accum2_acc_1827_nl = nl_Accum2_acc_1827_nl[9:0];
  assign nl_Product1_1_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[179:175]));
  assign Product1_1_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_590_nl = ({Accum2_acc_1827_nl , (Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_590_nl = nl_Accum2_acc_590_nl[15:0];
  assign nl_Accum2_acc_594_nl = Accum2_acc_591_nl + Accum2_acc_590_nl;
  assign Accum2_acc_594_nl = nl_Accum2_acc_594_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1 = Accum2_acc_595_nl
      + Accum2_acc_594_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[824:820]));
  assign Product1_2_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1464:1460]));
  assign Product1_3_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_602_nl = (readslicef_20_16_4(Product1_2_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_602_nl = nl_Accum2_acc_602_nl[15:0];
  assign nl_Product1_4_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2104:2100]));
  assign Product1_4_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2744:2740]));
  assign Product1_5_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_601_nl = (readslicef_20_16_4(Product1_4_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_601_nl = nl_Accum2_acc_601_nl[15:0];
  assign nl_Product1_6_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3384:3380]));
  assign Product1_6_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4024:4020]));
  assign Product1_7_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_600_nl = (readslicef_20_16_4(Product1_6_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_600_nl = nl_Accum2_acc_600_nl[15:0];
  assign nl_Product1_8_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4664:4660]));
  assign Product1_8_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5304:5300]));
  assign Product1_9_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_599_nl = (readslicef_20_16_4(Product1_8_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_599_nl = nl_Accum2_acc_599_nl[15:0];
  assign nl_Accum2_acc_608_nl = Accum2_acc_602_nl + Accum2_acc_601_nl + Accum2_acc_600_nl
      + Accum2_acc_599_nl;
  assign Accum2_acc_608_nl = nl_Accum2_acc_608_nl[15:0];
  assign nl_Product1_10_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5944:5940]));
  assign Product1_10_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6584:6580]));
  assign Product1_11_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_598_nl = (readslicef_20_16_4(Product1_10_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_598_nl = nl_Accum2_acc_598_nl[15:0];
  assign nl_Product1_12_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7224:7220]));
  assign Product1_12_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7864:7860]));
  assign Product1_13_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_597_nl = (readslicef_20_16_4(Product1_12_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_597_nl = nl_Accum2_acc_597_nl[15:0];
  assign nl_Accum2_acc_604_nl = Accum2_acc_598_nl + Accum2_acc_597_nl;
  assign Accum2_acc_604_nl = nl_Accum2_acc_604_nl[15:0];
  assign nl_Accum2_acc_1828_nl = (Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[184:180]);
  assign Accum2_acc_1828_nl = nl_Accum2_acc_1828_nl[9:0];
  assign nl_Product1_1_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[184:180]));
  assign Product1_1_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_603_nl = ({Accum2_acc_1828_nl , (Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_603_nl = nl_Accum2_acc_603_nl[15:0];
  assign nl_Accum2_acc_607_nl = Accum2_acc_604_nl + Accum2_acc_603_nl;
  assign Accum2_acc_607_nl = nl_Accum2_acc_607_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1 = Accum2_acc_608_nl
      + Accum2_acc_607_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[829:825]));
  assign Product1_2_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1469:1465]));
  assign Product1_3_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_615_nl = (readslicef_20_16_4(Product1_2_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_615_nl = nl_Accum2_acc_615_nl[15:0];
  assign nl_Product1_4_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2109:2105]));
  assign Product1_4_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2749:2745]));
  assign Product1_5_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_614_nl = (readslicef_20_16_4(Product1_4_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_614_nl = nl_Accum2_acc_614_nl[15:0];
  assign nl_Product1_6_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3389:3385]));
  assign Product1_6_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4029:4025]));
  assign Product1_7_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_613_nl = (readslicef_20_16_4(Product1_6_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_613_nl = nl_Accum2_acc_613_nl[15:0];
  assign nl_Product1_8_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4669:4665]));
  assign Product1_8_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5309:5305]));
  assign Product1_9_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_612_nl = (readslicef_20_16_4(Product1_8_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_612_nl = nl_Accum2_acc_612_nl[15:0];
  assign nl_Accum2_acc_621_nl = Accum2_acc_615_nl + Accum2_acc_614_nl + Accum2_acc_613_nl
      + Accum2_acc_612_nl;
  assign Accum2_acc_621_nl = nl_Accum2_acc_621_nl[15:0];
  assign nl_Product1_10_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5949:5945]));
  assign Product1_10_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6589:6585]));
  assign Product1_11_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_611_nl = (readslicef_20_16_4(Product1_10_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_611_nl = nl_Accum2_acc_611_nl[15:0];
  assign nl_Product1_12_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7229:7225]));
  assign Product1_12_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7869:7865]));
  assign Product1_13_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_610_nl = (readslicef_20_16_4(Product1_12_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_610_nl = nl_Accum2_acc_610_nl[15:0];
  assign nl_Accum2_acc_617_nl = Accum2_acc_611_nl + Accum2_acc_610_nl;
  assign Accum2_acc_617_nl = nl_Accum2_acc_617_nl[15:0];
  assign nl_Accum2_acc_1829_nl = (Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[189:185]);
  assign Accum2_acc_1829_nl = nl_Accum2_acc_1829_nl[9:0];
  assign nl_Product1_1_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[189:185]));
  assign Product1_1_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_616_nl = ({Accum2_acc_1829_nl , (Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_616_nl = nl_Accum2_acc_616_nl[15:0];
  assign nl_Accum2_acc_620_nl = Accum2_acc_617_nl + Accum2_acc_616_nl;
  assign Accum2_acc_620_nl = nl_Accum2_acc_620_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1 = Accum2_acc_621_nl
      + Accum2_acc_620_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[834:830]));
  assign Product1_2_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1474:1470]));
  assign Product1_3_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_628_nl = (readslicef_20_16_4(Product1_2_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_628_nl = nl_Accum2_acc_628_nl[15:0];
  assign nl_Product1_4_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2114:2110]));
  assign Product1_4_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2754:2750]));
  assign Product1_5_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_627_nl = (readslicef_20_16_4(Product1_4_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_627_nl = nl_Accum2_acc_627_nl[15:0];
  assign nl_Product1_6_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3394:3390]));
  assign Product1_6_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4034:4030]));
  assign Product1_7_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_626_nl = (readslicef_20_16_4(Product1_6_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_626_nl = nl_Accum2_acc_626_nl[15:0];
  assign nl_Product1_8_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4674:4670]));
  assign Product1_8_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5314:5310]));
  assign Product1_9_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_625_nl = (readslicef_20_16_4(Product1_8_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_625_nl = nl_Accum2_acc_625_nl[15:0];
  assign nl_Accum2_acc_634_nl = Accum2_acc_628_nl + Accum2_acc_627_nl + Accum2_acc_626_nl
      + Accum2_acc_625_nl;
  assign Accum2_acc_634_nl = nl_Accum2_acc_634_nl[15:0];
  assign nl_Product1_10_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5954:5950]));
  assign Product1_10_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6594:6590]));
  assign Product1_11_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_624_nl = (readslicef_20_16_4(Product1_10_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_624_nl = nl_Accum2_acc_624_nl[15:0];
  assign nl_Product1_12_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7234:7230]));
  assign Product1_12_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7874:7870]));
  assign Product1_13_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_623_nl = (readslicef_20_16_4(Product1_12_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_623_nl = nl_Accum2_acc_623_nl[15:0];
  assign nl_Accum2_acc_630_nl = Accum2_acc_624_nl + Accum2_acc_623_nl;
  assign Accum2_acc_630_nl = nl_Accum2_acc_630_nl[15:0];
  assign nl_Accum2_acc_1830_nl = (Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[194:190]);
  assign Accum2_acc_1830_nl = nl_Accum2_acc_1830_nl[9:0];
  assign nl_Product1_1_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[194:190]));
  assign Product1_1_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_629_nl = ({Accum2_acc_1830_nl , (Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_629_nl = nl_Accum2_acc_629_nl[15:0];
  assign nl_Accum2_acc_633_nl = Accum2_acc_630_nl + Accum2_acc_629_nl;
  assign Accum2_acc_633_nl = nl_Accum2_acc_633_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1 = Accum2_acc_634_nl
      + Accum2_acc_633_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[839:835]));
  assign Product1_2_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1479:1475]));
  assign Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_641_nl = (readslicef_20_16_4(Product1_2_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_641_nl = nl_Accum2_acc_641_nl[15:0];
  assign nl_Product1_4_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2119:2115]));
  assign Product1_4_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2759:2755]));
  assign Product1_5_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_640_nl = (readslicef_20_16_4(Product1_4_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_640_nl = nl_Accum2_acc_640_nl[15:0];
  assign nl_Product1_6_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3399:3395]));
  assign Product1_6_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4039:4035]));
  assign Product1_7_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_639_nl = (readslicef_20_16_4(Product1_6_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_639_nl = nl_Accum2_acc_639_nl[15:0];
  assign nl_Product1_8_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4679:4675]));
  assign Product1_8_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5319:5315]));
  assign Product1_9_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_638_nl = (readslicef_20_16_4(Product1_8_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_638_nl = nl_Accum2_acc_638_nl[15:0];
  assign nl_Accum2_acc_647_nl = Accum2_acc_641_nl + Accum2_acc_640_nl + Accum2_acc_639_nl
      + Accum2_acc_638_nl;
  assign Accum2_acc_647_nl = nl_Accum2_acc_647_nl[15:0];
  assign nl_Product1_10_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5959:5955]));
  assign Product1_10_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6599:6595]));
  assign Product1_11_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_637_nl = (readslicef_20_16_4(Product1_10_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_637_nl = nl_Accum2_acc_637_nl[15:0];
  assign nl_Product1_12_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7239:7235]));
  assign Product1_12_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7879:7875]));
  assign Product1_13_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_636_nl = (readslicef_20_16_4(Product1_12_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_636_nl = nl_Accum2_acc_636_nl[15:0];
  assign nl_Accum2_acc_643_nl = Accum2_acc_637_nl + Accum2_acc_636_nl;
  assign Accum2_acc_643_nl = nl_Accum2_acc_643_nl[15:0];
  assign nl_Accum2_acc_1831_nl = (Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[199:195]);
  assign Accum2_acc_1831_nl = nl_Accum2_acc_1831_nl[9:0];
  assign nl_Product1_1_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[199:195]));
  assign Product1_1_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_642_nl = ({Accum2_acc_1831_nl , (Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_642_nl = nl_Accum2_acc_642_nl[15:0];
  assign nl_Accum2_acc_646_nl = Accum2_acc_643_nl + Accum2_acc_642_nl;
  assign Accum2_acc_646_nl = nl_Accum2_acc_646_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1 = Accum2_acc_647_nl
      + Accum2_acc_646_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[844:840]));
  assign Product1_2_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1484:1480]));
  assign Product1_3_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_654_nl = (readslicef_20_16_4(Product1_2_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_654_nl = nl_Accum2_acc_654_nl[15:0];
  assign nl_Product1_4_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2124:2120]));
  assign Product1_4_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2764:2760]));
  assign Product1_5_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_653_nl = (readslicef_20_16_4(Product1_4_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_653_nl = nl_Accum2_acc_653_nl[15:0];
  assign nl_Product1_6_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3404:3400]));
  assign Product1_6_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4044:4040]));
  assign Product1_7_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_652_nl = (readslicef_20_16_4(Product1_6_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_652_nl = nl_Accum2_acc_652_nl[15:0];
  assign nl_Product1_8_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4684:4680]));
  assign Product1_8_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5324:5320]));
  assign Product1_9_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_651_nl = (readslicef_20_16_4(Product1_8_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_651_nl = nl_Accum2_acc_651_nl[15:0];
  assign nl_Accum2_acc_660_nl = Accum2_acc_654_nl + Accum2_acc_653_nl + Accum2_acc_652_nl
      + Accum2_acc_651_nl;
  assign Accum2_acc_660_nl = nl_Accum2_acc_660_nl[15:0];
  assign nl_Product1_10_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5964:5960]));
  assign Product1_10_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6604:6600]));
  assign Product1_11_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_650_nl = (readslicef_20_16_4(Product1_10_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_650_nl = nl_Accum2_acc_650_nl[15:0];
  assign nl_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7244:7240]));
  assign Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7884:7880]));
  assign Product1_13_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_649_nl = (readslicef_20_16_4(Product1_12_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_649_nl = nl_Accum2_acc_649_nl[15:0];
  assign nl_Accum2_acc_656_nl = Accum2_acc_650_nl + Accum2_acc_649_nl;
  assign Accum2_acc_656_nl = nl_Accum2_acc_656_nl[15:0];
  assign nl_Accum2_acc_1832_nl = (Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[204:200]);
  assign Accum2_acc_1832_nl = nl_Accum2_acc_1832_nl[9:0];
  assign nl_Product1_1_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[204:200]));
  assign Product1_1_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_655_nl = ({Accum2_acc_1832_nl , (Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_655_nl = nl_Accum2_acc_655_nl[15:0];
  assign nl_Accum2_acc_659_nl = Accum2_acc_656_nl + Accum2_acc_655_nl;
  assign Accum2_acc_659_nl = nl_Accum2_acc_659_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1 = Accum2_acc_660_nl
      + Accum2_acc_659_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[849:845]));
  assign Product1_2_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1489:1485]));
  assign Product1_3_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_667_nl = (readslicef_20_16_4(Product1_2_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_667_nl = nl_Accum2_acc_667_nl[15:0];
  assign nl_Product1_4_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2129:2125]));
  assign Product1_4_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2769:2765]));
  assign Product1_5_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_666_nl = (readslicef_20_16_4(Product1_4_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_666_nl = nl_Accum2_acc_666_nl[15:0];
  assign nl_Product1_6_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3409:3405]));
  assign Product1_6_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4049:4045]));
  assign Product1_7_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_665_nl = (readslicef_20_16_4(Product1_6_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_665_nl = nl_Accum2_acc_665_nl[15:0];
  assign nl_Product1_8_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4689:4685]));
  assign Product1_8_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5329:5325]));
  assign Product1_9_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_664_nl = (readslicef_20_16_4(Product1_8_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_664_nl = nl_Accum2_acc_664_nl[15:0];
  assign nl_Accum2_acc_673_nl = Accum2_acc_667_nl + Accum2_acc_666_nl + Accum2_acc_665_nl
      + Accum2_acc_664_nl;
  assign Accum2_acc_673_nl = nl_Accum2_acc_673_nl[15:0];
  assign nl_Product1_10_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5969:5965]));
  assign Product1_10_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6609:6605]));
  assign Product1_11_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_663_nl = (readslicef_20_16_4(Product1_10_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_663_nl = nl_Accum2_acc_663_nl[15:0];
  assign nl_Product1_12_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7249:7245]));
  assign Product1_12_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7889:7885]));
  assign Product1_13_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_662_nl = (readslicef_20_16_4(Product1_12_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_662_nl = nl_Accum2_acc_662_nl[15:0];
  assign nl_Accum2_acc_669_nl = Accum2_acc_663_nl + Accum2_acc_662_nl;
  assign Accum2_acc_669_nl = nl_Accum2_acc_669_nl[15:0];
  assign nl_Accum2_acc_1833_nl = (Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[209:205]);
  assign Accum2_acc_1833_nl = nl_Accum2_acc_1833_nl[9:0];
  assign nl_Product1_1_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[209:205]));
  assign Product1_1_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_668_nl = ({Accum2_acc_1833_nl , (Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_668_nl = nl_Accum2_acc_668_nl[15:0];
  assign nl_Accum2_acc_672_nl = Accum2_acc_669_nl + Accum2_acc_668_nl;
  assign Accum2_acc_672_nl = nl_Accum2_acc_672_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1 = Accum2_acc_673_nl
      + Accum2_acc_672_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[854:850]));
  assign Product1_2_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1494:1490]));
  assign Product1_3_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_680_nl = (readslicef_20_16_4(Product1_2_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_680_nl = nl_Accum2_acc_680_nl[15:0];
  assign nl_Product1_4_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2134:2130]));
  assign Product1_4_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2774:2770]));
  assign Product1_5_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_679_nl = (readslicef_20_16_4(Product1_4_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_679_nl = nl_Accum2_acc_679_nl[15:0];
  assign nl_Product1_6_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3414:3410]));
  assign Product1_6_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4054:4050]));
  assign Product1_7_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_678_nl = (readslicef_20_16_4(Product1_6_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_678_nl = nl_Accum2_acc_678_nl[15:0];
  assign nl_Product1_8_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4694:4690]));
  assign Product1_8_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5334:5330]));
  assign Product1_9_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_677_nl = (readslicef_20_16_4(Product1_8_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_677_nl = nl_Accum2_acc_677_nl[15:0];
  assign nl_Accum2_acc_686_nl = Accum2_acc_680_nl + Accum2_acc_679_nl + Accum2_acc_678_nl
      + Accum2_acc_677_nl;
  assign Accum2_acc_686_nl = nl_Accum2_acc_686_nl[15:0];
  assign nl_Product1_10_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5974:5970]));
  assign Product1_10_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6614:6610]));
  assign Product1_11_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_676_nl = (readslicef_20_16_4(Product1_10_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_676_nl = nl_Accum2_acc_676_nl[15:0];
  assign nl_Product1_12_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7254:7250]));
  assign Product1_12_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7894:7890]));
  assign Product1_13_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_675_nl = (readslicef_20_16_4(Product1_12_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_675_nl = nl_Accum2_acc_675_nl[15:0];
  assign nl_Accum2_acc_682_nl = Accum2_acc_676_nl + Accum2_acc_675_nl;
  assign Accum2_acc_682_nl = nl_Accum2_acc_682_nl[15:0];
  assign nl_Accum2_acc_1834_nl = (Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[214:210]);
  assign Accum2_acc_1834_nl = nl_Accum2_acc_1834_nl[9:0];
  assign nl_Product1_1_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[214:210]));
  assign Product1_1_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_681_nl = ({Accum2_acc_1834_nl , (Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_681_nl = nl_Accum2_acc_681_nl[15:0];
  assign nl_Accum2_acc_685_nl = Accum2_acc_682_nl + Accum2_acc_681_nl;
  assign Accum2_acc_685_nl = nl_Accum2_acc_685_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1 = Accum2_acc_686_nl
      + Accum2_acc_685_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[859:855]));
  assign Product1_2_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1499:1495]));
  assign Product1_3_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_693_nl = (readslicef_20_16_4(Product1_2_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_693_nl = nl_Accum2_acc_693_nl[15:0];
  assign nl_Product1_4_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2139:2135]));
  assign Product1_4_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2779:2775]));
  assign Product1_5_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_692_nl = (readslicef_20_16_4(Product1_4_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_692_nl = nl_Accum2_acc_692_nl[15:0];
  assign nl_Product1_6_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3419:3415]));
  assign Product1_6_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4059:4055]));
  assign Product1_7_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_691_nl = (readslicef_20_16_4(Product1_6_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_691_nl = nl_Accum2_acc_691_nl[15:0];
  assign nl_Product1_8_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4699:4695]));
  assign Product1_8_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5339:5335]));
  assign Product1_9_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_690_nl = (readslicef_20_16_4(Product1_8_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_690_nl = nl_Accum2_acc_690_nl[15:0];
  assign nl_Accum2_acc_699_nl = Accum2_acc_693_nl + Accum2_acc_692_nl + Accum2_acc_691_nl
      + Accum2_acc_690_nl;
  assign Accum2_acc_699_nl = nl_Accum2_acc_699_nl[15:0];
  assign nl_Product1_10_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5979:5975]));
  assign Product1_10_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6619:6615]));
  assign Product1_11_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_689_nl = (readslicef_20_16_4(Product1_10_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_689_nl = nl_Accum2_acc_689_nl[15:0];
  assign nl_Product1_12_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7259:7255]));
  assign Product1_12_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7899:7895]));
  assign Product1_13_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_688_nl = (readslicef_20_16_4(Product1_12_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_688_nl = nl_Accum2_acc_688_nl[15:0];
  assign nl_Accum2_acc_695_nl = Accum2_acc_689_nl + Accum2_acc_688_nl;
  assign Accum2_acc_695_nl = nl_Accum2_acc_695_nl[15:0];
  assign nl_Accum2_acc_1835_nl = (Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[219:215]);
  assign Accum2_acc_1835_nl = nl_Accum2_acc_1835_nl[9:0];
  assign nl_Product1_1_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[219:215]));
  assign Product1_1_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_694_nl = ({Accum2_acc_1835_nl , (Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_694_nl = nl_Accum2_acc_694_nl[15:0];
  assign nl_Accum2_acc_698_nl = Accum2_acc_695_nl + Accum2_acc_694_nl;
  assign Accum2_acc_698_nl = nl_Accum2_acc_698_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1 = Accum2_acc_699_nl
      + Accum2_acc_698_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[864:860]));
  assign Product1_2_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1504:1500]));
  assign Product1_3_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_706_nl = (readslicef_20_16_4(Product1_2_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_706_nl = nl_Accum2_acc_706_nl[15:0];
  assign nl_Product1_4_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2144:2140]));
  assign Product1_4_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2784:2780]));
  assign Product1_5_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_705_nl = (readslicef_20_16_4(Product1_4_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_705_nl = nl_Accum2_acc_705_nl[15:0];
  assign nl_Product1_6_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3424:3420]));
  assign Product1_6_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4064:4060]));
  assign Product1_7_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_704_nl = (readslicef_20_16_4(Product1_6_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_704_nl = nl_Accum2_acc_704_nl[15:0];
  assign nl_Product1_8_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4704:4700]));
  assign Product1_8_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5344:5340]));
  assign Product1_9_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_703_nl = (readslicef_20_16_4(Product1_8_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_703_nl = nl_Accum2_acc_703_nl[15:0];
  assign nl_Accum2_acc_712_nl = Accum2_acc_706_nl + Accum2_acc_705_nl + Accum2_acc_704_nl
      + Accum2_acc_703_nl;
  assign Accum2_acc_712_nl = nl_Accum2_acc_712_nl[15:0];
  assign nl_Product1_10_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5984:5980]));
  assign Product1_10_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6624:6620]));
  assign Product1_11_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_702_nl = (readslicef_20_16_4(Product1_10_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_702_nl = nl_Accum2_acc_702_nl[15:0];
  assign nl_Product1_12_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7264:7260]));
  assign Product1_12_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7904:7900]));
  assign Product1_13_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_701_nl = (readslicef_20_16_4(Product1_12_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_701_nl = nl_Accum2_acc_701_nl[15:0];
  assign nl_Accum2_acc_708_nl = Accum2_acc_702_nl + Accum2_acc_701_nl;
  assign Accum2_acc_708_nl = nl_Accum2_acc_708_nl[15:0];
  assign nl_Accum2_acc_1836_nl = (Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[224:220]);
  assign Accum2_acc_1836_nl = nl_Accum2_acc_1836_nl[9:0];
  assign nl_Product1_1_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[224:220]));
  assign Product1_1_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_707_nl = ({Accum2_acc_1836_nl , (Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_707_nl = nl_Accum2_acc_707_nl[15:0];
  assign nl_Accum2_acc_711_nl = Accum2_acc_708_nl + Accum2_acc_707_nl;
  assign Accum2_acc_711_nl = nl_Accum2_acc_711_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1 = Accum2_acc_712_nl
      + Accum2_acc_711_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[869:865]));
  assign Product1_2_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1509:1505]));
  assign Product1_3_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_719_nl = (readslicef_20_16_4(Product1_2_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_719_nl = nl_Accum2_acc_719_nl[15:0];
  assign nl_Product1_4_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2149:2145]));
  assign Product1_4_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2789:2785]));
  assign Product1_5_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_718_nl = (readslicef_20_16_4(Product1_4_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_718_nl = nl_Accum2_acc_718_nl[15:0];
  assign nl_Product1_6_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3429:3425]));
  assign Product1_6_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4069:4065]));
  assign Product1_7_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_717_nl = (readslicef_20_16_4(Product1_6_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_717_nl = nl_Accum2_acc_717_nl[15:0];
  assign nl_Product1_8_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4709:4705]));
  assign Product1_8_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5349:5345]));
  assign Product1_9_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_716_nl = (readslicef_20_16_4(Product1_8_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_716_nl = nl_Accum2_acc_716_nl[15:0];
  assign nl_Accum2_acc_725_nl = Accum2_acc_719_nl + Accum2_acc_718_nl + Accum2_acc_717_nl
      + Accum2_acc_716_nl;
  assign Accum2_acc_725_nl = nl_Accum2_acc_725_nl[15:0];
  assign nl_Product1_10_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5989:5985]));
  assign Product1_10_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6629:6625]));
  assign Product1_11_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_715_nl = (readslicef_20_16_4(Product1_10_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_715_nl = nl_Accum2_acc_715_nl[15:0];
  assign nl_Product1_12_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7269:7265]));
  assign Product1_12_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7909:7905]));
  assign Product1_13_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_714_nl = (readslicef_20_16_4(Product1_12_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_714_nl = nl_Accum2_acc_714_nl[15:0];
  assign nl_Accum2_acc_721_nl = Accum2_acc_715_nl + Accum2_acc_714_nl;
  assign Accum2_acc_721_nl = nl_Accum2_acc_721_nl[15:0];
  assign nl_Accum2_acc_1837_nl = (Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[229:225]);
  assign Accum2_acc_1837_nl = nl_Accum2_acc_1837_nl[9:0];
  assign nl_Product1_1_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[229:225]));
  assign Product1_1_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_720_nl = ({Accum2_acc_1837_nl , (Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_720_nl = nl_Accum2_acc_720_nl[15:0];
  assign nl_Accum2_acc_724_nl = Accum2_acc_721_nl + Accum2_acc_720_nl;
  assign Accum2_acc_724_nl = nl_Accum2_acc_724_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1 = Accum2_acc_725_nl
      + Accum2_acc_724_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[874:870]));
  assign Product1_2_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1514:1510]));
  assign Product1_3_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_732_nl = (readslicef_20_16_4(Product1_2_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_732_nl = nl_Accum2_acc_732_nl[15:0];
  assign nl_Product1_4_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2154:2150]));
  assign Product1_4_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2794:2790]));
  assign Product1_5_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_731_nl = (readslicef_20_16_4(Product1_4_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_731_nl = nl_Accum2_acc_731_nl[15:0];
  assign nl_Product1_6_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3434:3430]));
  assign Product1_6_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4074:4070]));
  assign Product1_7_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_730_nl = (readslicef_20_16_4(Product1_6_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_730_nl = nl_Accum2_acc_730_nl[15:0];
  assign nl_Product1_8_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4714:4710]));
  assign Product1_8_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5354:5350]));
  assign Product1_9_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_729_nl = (readslicef_20_16_4(Product1_8_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_729_nl = nl_Accum2_acc_729_nl[15:0];
  assign nl_Accum2_acc_738_nl = Accum2_acc_732_nl + Accum2_acc_731_nl + Accum2_acc_730_nl
      + Accum2_acc_729_nl;
  assign Accum2_acc_738_nl = nl_Accum2_acc_738_nl[15:0];
  assign nl_Product1_10_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5994:5990]));
  assign Product1_10_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6634:6630]));
  assign Product1_11_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_728_nl = (readslicef_20_16_4(Product1_10_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_728_nl = nl_Accum2_acc_728_nl[15:0];
  assign nl_Product1_12_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7274:7270]));
  assign Product1_12_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7914:7910]));
  assign Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_727_nl = (readslicef_20_16_4(Product1_12_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_727_nl = nl_Accum2_acc_727_nl[15:0];
  assign nl_Accum2_acc_734_nl = Accum2_acc_728_nl + Accum2_acc_727_nl;
  assign Accum2_acc_734_nl = nl_Accum2_acc_734_nl[15:0];
  assign nl_Accum2_acc_1838_nl = (Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[234:230]);
  assign Accum2_acc_1838_nl = nl_Accum2_acc_1838_nl[9:0];
  assign nl_Product1_1_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[234:230]));
  assign Product1_1_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_733_nl = ({Accum2_acc_1838_nl , (Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_733_nl = nl_Accum2_acc_733_nl[15:0];
  assign nl_Accum2_acc_737_nl = Accum2_acc_734_nl + Accum2_acc_733_nl;
  assign Accum2_acc_737_nl = nl_Accum2_acc_737_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1 = Accum2_acc_738_nl
      + Accum2_acc_737_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[879:875]));
  assign Product1_2_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1519:1515]));
  assign Product1_3_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_745_nl = (readslicef_20_16_4(Product1_2_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_745_nl = nl_Accum2_acc_745_nl[15:0];
  assign nl_Product1_4_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2159:2155]));
  assign Product1_4_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2799:2795]));
  assign Product1_5_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_744_nl = (readslicef_20_16_4(Product1_4_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_744_nl = nl_Accum2_acc_744_nl[15:0];
  assign nl_Product1_6_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3439:3435]));
  assign Product1_6_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4079:4075]));
  assign Product1_7_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_743_nl = (readslicef_20_16_4(Product1_6_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_743_nl = nl_Accum2_acc_743_nl[15:0];
  assign nl_Product1_8_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4719:4715]));
  assign Product1_8_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5359:5355]));
  assign Product1_9_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_742_nl = (readslicef_20_16_4(Product1_8_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_742_nl = nl_Accum2_acc_742_nl[15:0];
  assign nl_Accum2_acc_751_nl = Accum2_acc_745_nl + Accum2_acc_744_nl + Accum2_acc_743_nl
      + Accum2_acc_742_nl;
  assign Accum2_acc_751_nl = nl_Accum2_acc_751_nl[15:0];
  assign nl_Product1_10_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[5999:5995]));
  assign Product1_10_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6639:6635]));
  assign Product1_11_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_741_nl = (readslicef_20_16_4(Product1_10_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_741_nl = nl_Accum2_acc_741_nl[15:0];
  assign nl_Product1_12_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7279:7275]));
  assign Product1_12_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7919:7915]));
  assign Product1_13_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_740_nl = (readslicef_20_16_4(Product1_12_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_740_nl = nl_Accum2_acc_740_nl[15:0];
  assign nl_Accum2_acc_747_nl = Accum2_acc_741_nl + Accum2_acc_740_nl;
  assign Accum2_acc_747_nl = nl_Accum2_acc_747_nl[15:0];
  assign nl_Accum2_acc_1839_nl = (Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[239:235]);
  assign Accum2_acc_1839_nl = nl_Accum2_acc_1839_nl[9:0];
  assign nl_Product1_1_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[239:235]));
  assign Product1_1_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_746_nl = ({Accum2_acc_1839_nl , (Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_746_nl = nl_Accum2_acc_746_nl[15:0];
  assign nl_Accum2_acc_750_nl = Accum2_acc_747_nl + Accum2_acc_746_nl;
  assign Accum2_acc_750_nl = nl_Accum2_acc_750_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1 = Accum2_acc_751_nl
      + Accum2_acc_750_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[884:880]));
  assign Product1_2_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1524:1520]));
  assign Product1_3_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_758_nl = (readslicef_20_16_4(Product1_2_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_758_nl = nl_Accum2_acc_758_nl[15:0];
  assign nl_Product1_4_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2164:2160]));
  assign Product1_4_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2804:2800]));
  assign Product1_5_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_757_nl = (readslicef_20_16_4(Product1_4_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_757_nl = nl_Accum2_acc_757_nl[15:0];
  assign nl_Product1_6_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3444:3440]));
  assign Product1_6_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4084:4080]));
  assign Product1_7_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_756_nl = (readslicef_20_16_4(Product1_6_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_756_nl = nl_Accum2_acc_756_nl[15:0];
  assign nl_Product1_8_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4724:4720]));
  assign Product1_8_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5364:5360]));
  assign Product1_9_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_755_nl = (readslicef_20_16_4(Product1_8_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_755_nl = nl_Accum2_acc_755_nl[15:0];
  assign nl_Accum2_acc_764_nl = Accum2_acc_758_nl + Accum2_acc_757_nl + Accum2_acc_756_nl
      + Accum2_acc_755_nl;
  assign Accum2_acc_764_nl = nl_Accum2_acc_764_nl[15:0];
  assign nl_Product1_10_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6004:6000]));
  assign Product1_10_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6644:6640]));
  assign Product1_11_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_754_nl = (readslicef_20_16_4(Product1_10_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_754_nl = nl_Accum2_acc_754_nl[15:0];
  assign nl_Product1_12_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7284:7280]));
  assign Product1_12_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7924:7920]));
  assign Product1_13_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_753_nl = (readslicef_20_16_4(Product1_12_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_753_nl = nl_Accum2_acc_753_nl[15:0];
  assign nl_Accum2_acc_760_nl = Accum2_acc_754_nl + Accum2_acc_753_nl;
  assign Accum2_acc_760_nl = nl_Accum2_acc_760_nl[15:0];
  assign nl_Accum2_acc_1840_nl = (Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[244:240]);
  assign Accum2_acc_1840_nl = nl_Accum2_acc_1840_nl[9:0];
  assign nl_Product1_1_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[244:240]));
  assign Product1_1_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_759_nl = ({Accum2_acc_1840_nl , (Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_759_nl = nl_Accum2_acc_759_nl[15:0];
  assign nl_Accum2_acc_763_nl = Accum2_acc_760_nl + Accum2_acc_759_nl;
  assign Accum2_acc_763_nl = nl_Accum2_acc_763_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1 = Accum2_acc_764_nl
      + Accum2_acc_763_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[889:885]));
  assign Product1_2_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1529:1525]));
  assign Product1_3_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_771_nl = (readslicef_20_16_4(Product1_2_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_771_nl = nl_Accum2_acc_771_nl[15:0];
  assign nl_Product1_4_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2169:2165]));
  assign Product1_4_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2809:2805]));
  assign Product1_5_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_770_nl = (readslicef_20_16_4(Product1_4_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_770_nl = nl_Accum2_acc_770_nl[15:0];
  assign nl_Product1_6_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3449:3445]));
  assign Product1_6_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4089:4085]));
  assign Product1_7_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_769_nl = (readslicef_20_16_4(Product1_6_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_769_nl = nl_Accum2_acc_769_nl[15:0];
  assign nl_Product1_8_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4729:4725]));
  assign Product1_8_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5369:5365]));
  assign Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_768_nl = (readslicef_20_16_4(Product1_8_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_768_nl = nl_Accum2_acc_768_nl[15:0];
  assign nl_Accum2_acc_777_nl = Accum2_acc_771_nl + Accum2_acc_770_nl + Accum2_acc_769_nl
      + Accum2_acc_768_nl;
  assign Accum2_acc_777_nl = nl_Accum2_acc_777_nl[15:0];
  assign nl_Product1_10_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6009:6005]));
  assign Product1_10_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6649:6645]));
  assign Product1_11_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_767_nl = (readslicef_20_16_4(Product1_10_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_767_nl = nl_Accum2_acc_767_nl[15:0];
  assign nl_Product1_12_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7289:7285]));
  assign Product1_12_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7929:7925]));
  assign Product1_13_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_766_nl = (readslicef_20_16_4(Product1_12_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_766_nl = nl_Accum2_acc_766_nl[15:0];
  assign nl_Accum2_acc_773_nl = Accum2_acc_767_nl + Accum2_acc_766_nl;
  assign Accum2_acc_773_nl = nl_Accum2_acc_773_nl[15:0];
  assign nl_Accum2_acc_1841_nl = (Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[249:245]);
  assign Accum2_acc_1841_nl = nl_Accum2_acc_1841_nl[9:0];
  assign nl_Product1_1_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[249:245]));
  assign Product1_1_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_772_nl = ({Accum2_acc_1841_nl , (Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_772_nl = nl_Accum2_acc_772_nl[15:0];
  assign nl_Accum2_acc_776_nl = Accum2_acc_773_nl + Accum2_acc_772_nl;
  assign Accum2_acc_776_nl = nl_Accum2_acc_776_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1 = Accum2_acc_777_nl
      + Accum2_acc_776_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[894:890]));
  assign Product1_2_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1534:1530]));
  assign Product1_3_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_784_nl = (readslicef_20_16_4(Product1_2_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_784_nl = nl_Accum2_acc_784_nl[15:0];
  assign nl_Product1_4_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2174:2170]));
  assign Product1_4_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2814:2810]));
  assign Product1_5_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_783_nl = (readslicef_20_16_4(Product1_4_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_783_nl = nl_Accum2_acc_783_nl[15:0];
  assign nl_Product1_6_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3454:3450]));
  assign Product1_6_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4094:4090]));
  assign Product1_7_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_782_nl = (readslicef_20_16_4(Product1_6_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_782_nl = nl_Accum2_acc_782_nl[15:0];
  assign nl_Product1_8_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4734:4730]));
  assign Product1_8_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5374:5370]));
  assign Product1_9_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_781_nl = (readslicef_20_16_4(Product1_8_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_781_nl = nl_Accum2_acc_781_nl[15:0];
  assign nl_Accum2_acc_790_nl = Accum2_acc_784_nl + Accum2_acc_783_nl + Accum2_acc_782_nl
      + Accum2_acc_781_nl;
  assign Accum2_acc_790_nl = nl_Accum2_acc_790_nl[15:0];
  assign nl_Product1_10_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6014:6010]));
  assign Product1_10_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6654:6650]));
  assign Product1_11_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_780_nl = (readslicef_20_16_4(Product1_10_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_780_nl = nl_Accum2_acc_780_nl[15:0];
  assign nl_Product1_12_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7294:7290]));
  assign Product1_12_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7934:7930]));
  assign Product1_13_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_779_nl = (readslicef_20_16_4(Product1_12_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_779_nl = nl_Accum2_acc_779_nl[15:0];
  assign nl_Accum2_acc_786_nl = Accum2_acc_780_nl + Accum2_acc_779_nl;
  assign Accum2_acc_786_nl = nl_Accum2_acc_786_nl[15:0];
  assign nl_Accum2_acc_1842_nl = (Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[254:250]);
  assign Accum2_acc_1842_nl = nl_Accum2_acc_1842_nl[9:0];
  assign nl_Product1_1_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[254:250]));
  assign Product1_1_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_785_nl = ({Accum2_acc_1842_nl , (Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_785_nl = nl_Accum2_acc_785_nl[15:0];
  assign nl_Accum2_acc_789_nl = Accum2_acc_786_nl + Accum2_acc_785_nl;
  assign Accum2_acc_789_nl = nl_Accum2_acc_789_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1 = Accum2_acc_790_nl
      + Accum2_acc_789_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[899:895]));
  assign Product1_2_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1539:1535]));
  assign Product1_3_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_797_nl = (readslicef_20_16_4(Product1_2_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_797_nl = nl_Accum2_acc_797_nl[15:0];
  assign nl_Product1_4_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2179:2175]));
  assign Product1_4_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2819:2815]));
  assign Product1_5_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_796_nl = (readslicef_20_16_4(Product1_4_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_796_nl = nl_Accum2_acc_796_nl[15:0];
  assign nl_Product1_6_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3459:3455]));
  assign Product1_6_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4099:4095]));
  assign Product1_7_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_795_nl = (readslicef_20_16_4(Product1_6_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_795_nl = nl_Accum2_acc_795_nl[15:0];
  assign nl_Product1_8_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4739:4735]));
  assign Product1_8_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5379:5375]));
  assign Product1_9_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_794_nl = (readslicef_20_16_4(Product1_8_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_794_nl = nl_Accum2_acc_794_nl[15:0];
  assign nl_Accum2_acc_803_nl = Accum2_acc_797_nl + Accum2_acc_796_nl + Accum2_acc_795_nl
      + Accum2_acc_794_nl;
  assign Accum2_acc_803_nl = nl_Accum2_acc_803_nl[15:0];
  assign nl_Product1_10_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6019:6015]));
  assign Product1_10_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6659:6655]));
  assign Product1_11_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_793_nl = (readslicef_20_16_4(Product1_10_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_793_nl = nl_Accum2_acc_793_nl[15:0];
  assign nl_Product1_12_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7299:7295]));
  assign Product1_12_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7939:7935]));
  assign Product1_13_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_792_nl = (readslicef_20_16_4(Product1_12_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_792_nl = nl_Accum2_acc_792_nl[15:0];
  assign nl_Accum2_acc_799_nl = Accum2_acc_793_nl + Accum2_acc_792_nl;
  assign Accum2_acc_799_nl = nl_Accum2_acc_799_nl[15:0];
  assign nl_Accum2_acc_1843_nl = (Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[259:255]);
  assign Accum2_acc_1843_nl = nl_Accum2_acc_1843_nl[9:0];
  assign nl_Product1_1_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[259:255]));
  assign Product1_1_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_798_nl = ({Accum2_acc_1843_nl , (Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_798_nl = nl_Accum2_acc_798_nl[15:0];
  assign nl_Accum2_acc_802_nl = Accum2_acc_799_nl + Accum2_acc_798_nl;
  assign Accum2_acc_802_nl = nl_Accum2_acc_802_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1 = Accum2_acc_803_nl
      + Accum2_acc_802_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[904:900]));
  assign Product1_2_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1544:1540]));
  assign Product1_3_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_810_nl = (readslicef_20_16_4(Product1_2_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_810_nl = nl_Accum2_acc_810_nl[15:0];
  assign nl_Product1_4_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2184:2180]));
  assign Product1_4_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2824:2820]));
  assign Product1_5_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_809_nl = (readslicef_20_16_4(Product1_4_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_809_nl = nl_Accum2_acc_809_nl[15:0];
  assign nl_Product1_6_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3464:3460]));
  assign Product1_6_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4104:4100]));
  assign Product1_7_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_808_nl = (readslicef_20_16_4(Product1_6_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_808_nl = nl_Accum2_acc_808_nl[15:0];
  assign nl_Product1_8_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4744:4740]));
  assign Product1_8_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5384:5380]));
  assign Product1_9_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_807_nl = (readslicef_20_16_4(Product1_8_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_807_nl = nl_Accum2_acc_807_nl[15:0];
  assign nl_Accum2_acc_816_nl = Accum2_acc_810_nl + Accum2_acc_809_nl + Accum2_acc_808_nl
      + Accum2_acc_807_nl;
  assign Accum2_acc_816_nl = nl_Accum2_acc_816_nl[15:0];
  assign nl_Product1_10_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6024:6020]));
  assign Product1_10_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6664:6660]));
  assign Product1_11_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_806_nl = (readslicef_20_16_4(Product1_10_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_806_nl = nl_Accum2_acc_806_nl[15:0];
  assign nl_Product1_12_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7304:7300]));
  assign Product1_12_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7944:7940]));
  assign Product1_13_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_805_nl = (readslicef_20_16_4(Product1_12_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_805_nl = nl_Accum2_acc_805_nl[15:0];
  assign nl_Accum2_acc_812_nl = Accum2_acc_806_nl + Accum2_acc_805_nl;
  assign Accum2_acc_812_nl = nl_Accum2_acc_812_nl[15:0];
  assign nl_Accum2_acc_1844_nl = (Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[264:260]);
  assign Accum2_acc_1844_nl = nl_Accum2_acc_1844_nl[9:0];
  assign nl_Product1_1_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[264:260]));
  assign Product1_1_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_811_nl = ({Accum2_acc_1844_nl , (Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_811_nl = nl_Accum2_acc_811_nl[15:0];
  assign nl_Accum2_acc_815_nl = Accum2_acc_812_nl + Accum2_acc_811_nl;
  assign Accum2_acc_815_nl = nl_Accum2_acc_815_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1 = Accum2_acc_816_nl
      + Accum2_acc_815_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[909:905]));
  assign Product1_2_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1549:1545]));
  assign Product1_3_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_823_nl = (readslicef_20_16_4(Product1_2_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_823_nl = nl_Accum2_acc_823_nl[15:0];
  assign nl_Product1_4_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2189:2185]));
  assign Product1_4_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2829:2825]));
  assign Product1_5_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_822_nl = (readslicef_20_16_4(Product1_4_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_822_nl = nl_Accum2_acc_822_nl[15:0];
  assign nl_Product1_6_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3469:3465]));
  assign Product1_6_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4109:4105]));
  assign Product1_7_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_821_nl = (readslicef_20_16_4(Product1_6_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_821_nl = nl_Accum2_acc_821_nl[15:0];
  assign nl_Product1_8_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4749:4745]));
  assign Product1_8_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5389:5385]));
  assign Product1_9_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_820_nl = (readslicef_20_16_4(Product1_8_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_820_nl = nl_Accum2_acc_820_nl[15:0];
  assign nl_Accum2_acc_829_nl = Accum2_acc_823_nl + Accum2_acc_822_nl + Accum2_acc_821_nl
      + Accum2_acc_820_nl;
  assign Accum2_acc_829_nl = nl_Accum2_acc_829_nl[15:0];
  assign nl_Product1_10_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6029:6025]));
  assign Product1_10_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6669:6665]));
  assign Product1_11_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_819_nl = (readslicef_20_16_4(Product1_10_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_819_nl = nl_Accum2_acc_819_nl[15:0];
  assign nl_Product1_12_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7309:7305]));
  assign Product1_12_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7949:7945]));
  assign Product1_13_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_818_nl = (readslicef_20_16_4(Product1_12_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_818_nl = nl_Accum2_acc_818_nl[15:0];
  assign nl_Accum2_acc_825_nl = Accum2_acc_819_nl + Accum2_acc_818_nl;
  assign Accum2_acc_825_nl = nl_Accum2_acc_825_nl[15:0];
  assign nl_Accum2_acc_1845_nl = (Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[269:265]);
  assign Accum2_acc_1845_nl = nl_Accum2_acc_1845_nl[9:0];
  assign nl_Product1_1_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[269:265]));
  assign Product1_1_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_824_nl = ({Accum2_acc_1845_nl , (Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_824_nl = nl_Accum2_acc_824_nl[15:0];
  assign nl_Accum2_acc_828_nl = Accum2_acc_825_nl + Accum2_acc_824_nl;
  assign Accum2_acc_828_nl = nl_Accum2_acc_828_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1 = Accum2_acc_829_nl
      + Accum2_acc_828_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[914:910]));
  assign Product1_2_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1554:1550]));
  assign Product1_3_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_836_nl = (readslicef_20_16_4(Product1_2_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_836_nl = nl_Accum2_acc_836_nl[15:0];
  assign nl_Product1_4_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2194:2190]));
  assign Product1_4_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2834:2830]));
  assign Product1_5_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_835_nl = (readslicef_20_16_4(Product1_4_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_835_nl = nl_Accum2_acc_835_nl[15:0];
  assign nl_Product1_6_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3474:3470]));
  assign Product1_6_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4114:4110]));
  assign Product1_7_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_834_nl = (readslicef_20_16_4(Product1_6_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_834_nl = nl_Accum2_acc_834_nl[15:0];
  assign nl_Product1_8_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4754:4750]));
  assign Product1_8_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5394:5390]));
  assign Product1_9_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_833_nl = (readslicef_20_16_4(Product1_8_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_833_nl = nl_Accum2_acc_833_nl[15:0];
  assign nl_Accum2_acc_842_nl = Accum2_acc_836_nl + Accum2_acc_835_nl + Accum2_acc_834_nl
      + Accum2_acc_833_nl;
  assign Accum2_acc_842_nl = nl_Accum2_acc_842_nl[15:0];
  assign nl_Product1_10_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6034:6030]));
  assign Product1_10_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6674:6670]));
  assign Product1_11_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_832_nl = (readslicef_20_16_4(Product1_10_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_832_nl = nl_Accum2_acc_832_nl[15:0];
  assign nl_Product1_12_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7314:7310]));
  assign Product1_12_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7954:7950]));
  assign Product1_13_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_831_nl = (readslicef_20_16_4(Product1_12_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_831_nl = nl_Accum2_acc_831_nl[15:0];
  assign nl_Accum2_acc_838_nl = Accum2_acc_832_nl + Accum2_acc_831_nl;
  assign Accum2_acc_838_nl = nl_Accum2_acc_838_nl[15:0];
  assign nl_Accum2_acc_1846_nl = (Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[274:270]);
  assign Accum2_acc_1846_nl = nl_Accum2_acc_1846_nl[9:0];
  assign nl_Product1_1_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[274:270]));
  assign Product1_1_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_837_nl = ({Accum2_acc_1846_nl , (Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_837_nl = nl_Accum2_acc_837_nl[15:0];
  assign nl_Accum2_acc_841_nl = Accum2_acc_838_nl + Accum2_acc_837_nl;
  assign Accum2_acc_841_nl = nl_Accum2_acc_841_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1 = Accum2_acc_842_nl
      + Accum2_acc_841_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[919:915]));
  assign Product1_2_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1559:1555]));
  assign Product1_3_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_849_nl = (readslicef_20_16_4(Product1_2_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_849_nl = nl_Accum2_acc_849_nl[15:0];
  assign nl_Product1_4_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2199:2195]));
  assign Product1_4_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2839:2835]));
  assign Product1_5_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_848_nl = (readslicef_20_16_4(Product1_4_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_848_nl = nl_Accum2_acc_848_nl[15:0];
  assign nl_Product1_6_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3479:3475]));
  assign Product1_6_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4119:4115]));
  assign Product1_7_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_847_nl = (readslicef_20_16_4(Product1_6_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_847_nl = nl_Accum2_acc_847_nl[15:0];
  assign nl_Product1_8_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4759:4755]));
  assign Product1_8_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5399:5395]));
  assign Product1_9_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_846_nl = (readslicef_20_16_4(Product1_8_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_846_nl = nl_Accum2_acc_846_nl[15:0];
  assign nl_Accum2_acc_855_nl = Accum2_acc_849_nl + Accum2_acc_848_nl + Accum2_acc_847_nl
      + Accum2_acc_846_nl;
  assign Accum2_acc_855_nl = nl_Accum2_acc_855_nl[15:0];
  assign nl_Product1_10_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6039:6035]));
  assign Product1_10_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6679:6675]));
  assign Product1_11_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_845_nl = (readslicef_20_16_4(Product1_10_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_845_nl = nl_Accum2_acc_845_nl[15:0];
  assign nl_Product1_12_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7319:7315]));
  assign Product1_12_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7959:7955]));
  assign Product1_13_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_844_nl = (readslicef_20_16_4(Product1_12_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_844_nl = nl_Accum2_acc_844_nl[15:0];
  assign nl_Accum2_acc_851_nl = Accum2_acc_845_nl + Accum2_acc_844_nl;
  assign Accum2_acc_851_nl = nl_Accum2_acc_851_nl[15:0];
  assign nl_Accum2_acc_1847_nl = (Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[279:275]);
  assign Accum2_acc_1847_nl = nl_Accum2_acc_1847_nl[9:0];
  assign nl_Product1_1_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[279:275]));
  assign Product1_1_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_850_nl = ({Accum2_acc_1847_nl , (Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_850_nl = nl_Accum2_acc_850_nl[15:0];
  assign nl_Accum2_acc_854_nl = Accum2_acc_851_nl + Accum2_acc_850_nl;
  assign Accum2_acc_854_nl = nl_Accum2_acc_854_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1 = Accum2_acc_855_nl
      + Accum2_acc_854_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[924:920]));
  assign Product1_2_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1564:1560]));
  assign Product1_3_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_862_nl = (readslicef_20_16_4(Product1_2_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_862_nl = nl_Accum2_acc_862_nl[15:0];
  assign nl_Product1_4_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2204:2200]));
  assign Product1_4_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2844:2840]));
  assign Product1_5_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_861_nl = (readslicef_20_16_4(Product1_4_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_861_nl = nl_Accum2_acc_861_nl[15:0];
  assign nl_Product1_6_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3484:3480]));
  assign Product1_6_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4124:4120]));
  assign Product1_7_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_860_nl = (readslicef_20_16_4(Product1_6_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_860_nl = nl_Accum2_acc_860_nl[15:0];
  assign nl_Product1_8_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4764:4760]));
  assign Product1_8_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5404:5400]));
  assign Product1_9_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_859_nl = (readslicef_20_16_4(Product1_8_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_859_nl = nl_Accum2_acc_859_nl[15:0];
  assign nl_Accum2_acc_868_nl = Accum2_acc_862_nl + Accum2_acc_861_nl + Accum2_acc_860_nl
      + Accum2_acc_859_nl;
  assign Accum2_acc_868_nl = nl_Accum2_acc_868_nl[15:0];
  assign nl_Product1_10_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6044:6040]));
  assign Product1_10_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6684:6680]));
  assign Product1_11_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_858_nl = (readslicef_20_16_4(Product1_10_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_858_nl = nl_Accum2_acc_858_nl[15:0];
  assign nl_Product1_12_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7324:7320]));
  assign Product1_12_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7964:7960]));
  assign Product1_13_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_857_nl = (readslicef_20_16_4(Product1_12_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_857_nl = nl_Accum2_acc_857_nl[15:0];
  assign nl_Accum2_acc_864_nl = Accum2_acc_858_nl + Accum2_acc_857_nl;
  assign Accum2_acc_864_nl = nl_Accum2_acc_864_nl[15:0];
  assign nl_Accum2_acc_1848_nl = (Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[284:280]);
  assign Accum2_acc_1848_nl = nl_Accum2_acc_1848_nl[9:0];
  assign nl_Product1_1_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[284:280]));
  assign Product1_1_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_863_nl = ({Accum2_acc_1848_nl , (Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_863_nl = nl_Accum2_acc_863_nl[15:0];
  assign nl_Accum2_acc_867_nl = Accum2_acc_864_nl + Accum2_acc_863_nl;
  assign Accum2_acc_867_nl = nl_Accum2_acc_867_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1 = Accum2_acc_868_nl
      + Accum2_acc_867_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[929:925]));
  assign Product1_2_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1569:1565]));
  assign Product1_3_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_875_nl = (readslicef_20_16_4(Product1_2_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_875_nl = nl_Accum2_acc_875_nl[15:0];
  assign nl_Product1_4_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2209:2205]));
  assign Product1_4_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2849:2845]));
  assign Product1_5_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_874_nl = (readslicef_20_16_4(Product1_4_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_874_nl = nl_Accum2_acc_874_nl[15:0];
  assign nl_Product1_6_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3489:3485]));
  assign Product1_6_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4129:4125]));
  assign Product1_7_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_873_nl = (readslicef_20_16_4(Product1_6_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_873_nl = nl_Accum2_acc_873_nl[15:0];
  assign nl_Product1_8_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4769:4765]));
  assign Product1_8_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5409:5405]));
  assign Product1_9_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_872_nl = (readslicef_20_16_4(Product1_8_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_872_nl = nl_Accum2_acc_872_nl[15:0];
  assign nl_Accum2_acc_881_nl = Accum2_acc_875_nl + Accum2_acc_874_nl + Accum2_acc_873_nl
      + Accum2_acc_872_nl;
  assign Accum2_acc_881_nl = nl_Accum2_acc_881_nl[15:0];
  assign nl_Product1_10_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6049:6045]));
  assign Product1_10_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6689:6685]));
  assign Product1_11_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_871_nl = (readslicef_20_16_4(Product1_10_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_871_nl = nl_Accum2_acc_871_nl[15:0];
  assign nl_Product1_12_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7329:7325]));
  assign Product1_12_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7969:7965]));
  assign Product1_13_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_870_nl = (readslicef_20_16_4(Product1_12_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_870_nl = nl_Accum2_acc_870_nl[15:0];
  assign nl_Accum2_acc_877_nl = Accum2_acc_871_nl + Accum2_acc_870_nl;
  assign Accum2_acc_877_nl = nl_Accum2_acc_877_nl[15:0];
  assign nl_Accum2_acc_1849_nl = (Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[289:285]);
  assign Accum2_acc_1849_nl = nl_Accum2_acc_1849_nl[9:0];
  assign nl_Product1_1_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[289:285]));
  assign Product1_1_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_876_nl = ({Accum2_acc_1849_nl , (Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_876_nl = nl_Accum2_acc_876_nl[15:0];
  assign nl_Accum2_acc_880_nl = Accum2_acc_877_nl + Accum2_acc_876_nl;
  assign Accum2_acc_880_nl = nl_Accum2_acc_880_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1 = Accum2_acc_881_nl
      + Accum2_acc_880_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[934:930]));
  assign Product1_2_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1574:1570]));
  assign Product1_3_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_888_nl = (readslicef_20_16_4(Product1_2_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_888_nl = nl_Accum2_acc_888_nl[15:0];
  assign nl_Product1_4_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2214:2210]));
  assign Product1_4_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2854:2850]));
  assign Product1_5_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_887_nl = (readslicef_20_16_4(Product1_4_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_887_nl = nl_Accum2_acc_887_nl[15:0];
  assign nl_Product1_6_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3494:3490]));
  assign Product1_6_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4134:4130]));
  assign Product1_7_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_886_nl = (readslicef_20_16_4(Product1_6_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_886_nl = nl_Accum2_acc_886_nl[15:0];
  assign nl_Product1_8_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4774:4770]));
  assign Product1_8_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5414:5410]));
  assign Product1_9_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_885_nl = (readslicef_20_16_4(Product1_8_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_885_nl = nl_Accum2_acc_885_nl[15:0];
  assign nl_Accum2_acc_894_nl = Accum2_acc_888_nl + Accum2_acc_887_nl + Accum2_acc_886_nl
      + Accum2_acc_885_nl;
  assign Accum2_acc_894_nl = nl_Accum2_acc_894_nl[15:0];
  assign nl_Product1_10_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6054:6050]));
  assign Product1_10_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6694:6690]));
  assign Product1_11_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_884_nl = (readslicef_20_16_4(Product1_10_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_884_nl = nl_Accum2_acc_884_nl[15:0];
  assign nl_Product1_12_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7334:7330]));
  assign Product1_12_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7974:7970]));
  assign Product1_13_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_883_nl = (readslicef_20_16_4(Product1_12_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_883_nl = nl_Accum2_acc_883_nl[15:0];
  assign nl_Accum2_acc_890_nl = Accum2_acc_884_nl + Accum2_acc_883_nl;
  assign Accum2_acc_890_nl = nl_Accum2_acc_890_nl[15:0];
  assign nl_Accum2_acc_1850_nl = (Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[294:290]);
  assign Accum2_acc_1850_nl = nl_Accum2_acc_1850_nl[9:0];
  assign nl_Product1_1_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[294:290]));
  assign Product1_1_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_889_nl = ({Accum2_acc_1850_nl , (Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_889_nl = nl_Accum2_acc_889_nl[15:0];
  assign nl_Accum2_acc_893_nl = Accum2_acc_890_nl + Accum2_acc_889_nl;
  assign Accum2_acc_893_nl = nl_Accum2_acc_893_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1 = Accum2_acc_894_nl
      + Accum2_acc_893_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[939:935]));
  assign Product1_2_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1579:1575]));
  assign Product1_3_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_901_nl = (readslicef_20_16_4(Product1_2_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_901_nl = nl_Accum2_acc_901_nl[15:0];
  assign nl_Product1_4_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2219:2215]));
  assign Product1_4_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2859:2855]));
  assign Product1_5_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_900_nl = (readslicef_20_16_4(Product1_4_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_900_nl = nl_Accum2_acc_900_nl[15:0];
  assign nl_Product1_6_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3499:3495]));
  assign Product1_6_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4139:4135]));
  assign Product1_7_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_899_nl = (readslicef_20_16_4(Product1_6_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_899_nl = nl_Accum2_acc_899_nl[15:0];
  assign nl_Product1_8_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4779:4775]));
  assign Product1_8_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5419:5415]));
  assign Product1_9_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_898_nl = (readslicef_20_16_4(Product1_8_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_898_nl = nl_Accum2_acc_898_nl[15:0];
  assign nl_Accum2_acc_907_nl = Accum2_acc_901_nl + Accum2_acc_900_nl + Accum2_acc_899_nl
      + Accum2_acc_898_nl;
  assign Accum2_acc_907_nl = nl_Accum2_acc_907_nl[15:0];
  assign nl_Product1_10_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6059:6055]));
  assign Product1_10_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6699:6695]));
  assign Product1_11_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_897_nl = (readslicef_20_16_4(Product1_10_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_897_nl = nl_Accum2_acc_897_nl[15:0];
  assign nl_Product1_12_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7339:7335]));
  assign Product1_12_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7979:7975]));
  assign Product1_13_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_896_nl = (readslicef_20_16_4(Product1_12_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_896_nl = nl_Accum2_acc_896_nl[15:0];
  assign nl_Accum2_acc_903_nl = Accum2_acc_897_nl + Accum2_acc_896_nl;
  assign Accum2_acc_903_nl = nl_Accum2_acc_903_nl[15:0];
  assign nl_Accum2_acc_1851_nl = (Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[299:295]);
  assign Accum2_acc_1851_nl = nl_Accum2_acc_1851_nl[9:0];
  assign nl_Product1_1_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[299:295]));
  assign Product1_1_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_902_nl = ({Accum2_acc_1851_nl , (Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_902_nl = nl_Accum2_acc_902_nl[15:0];
  assign nl_Accum2_acc_906_nl = Accum2_acc_903_nl + Accum2_acc_902_nl;
  assign Accum2_acc_906_nl = nl_Accum2_acc_906_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1 = Accum2_acc_907_nl
      + Accum2_acc_906_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[944:940]));
  assign Product1_2_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1584:1580]));
  assign Product1_3_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_914_nl = (readslicef_20_16_4(Product1_2_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_914_nl = nl_Accum2_acc_914_nl[15:0];
  assign nl_Product1_4_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2224:2220]));
  assign Product1_4_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2864:2860]));
  assign Product1_5_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_913_nl = (readslicef_20_16_4(Product1_4_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_913_nl = nl_Accum2_acc_913_nl[15:0];
  assign nl_Product1_6_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3504:3500]));
  assign Product1_6_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4144:4140]));
  assign Product1_7_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_912_nl = (readslicef_20_16_4(Product1_6_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_912_nl = nl_Accum2_acc_912_nl[15:0];
  assign nl_Product1_8_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4784:4780]));
  assign Product1_8_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5424:5420]));
  assign Product1_9_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_911_nl = (readslicef_20_16_4(Product1_8_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_911_nl = nl_Accum2_acc_911_nl[15:0];
  assign nl_Accum2_acc_920_nl = Accum2_acc_914_nl + Accum2_acc_913_nl + Accum2_acc_912_nl
      + Accum2_acc_911_nl;
  assign Accum2_acc_920_nl = nl_Accum2_acc_920_nl[15:0];
  assign nl_Product1_10_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6064:6060]));
  assign Product1_10_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6704:6700]));
  assign Product1_11_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_910_nl = (readslicef_20_16_4(Product1_10_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_910_nl = nl_Accum2_acc_910_nl[15:0];
  assign nl_Product1_12_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7344:7340]));
  assign Product1_12_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7984:7980]));
  assign Product1_13_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_909_nl = (readslicef_20_16_4(Product1_12_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_909_nl = nl_Accum2_acc_909_nl[15:0];
  assign nl_Accum2_acc_916_nl = Accum2_acc_910_nl + Accum2_acc_909_nl;
  assign Accum2_acc_916_nl = nl_Accum2_acc_916_nl[15:0];
  assign nl_Accum2_acc_1852_nl = (Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[304:300]);
  assign Accum2_acc_1852_nl = nl_Accum2_acc_1852_nl[9:0];
  assign nl_Product1_1_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[304:300]));
  assign Product1_1_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_915_nl = ({Accum2_acc_1852_nl , (Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_915_nl = nl_Accum2_acc_915_nl[15:0];
  assign nl_Accum2_acc_919_nl = Accum2_acc_916_nl + Accum2_acc_915_nl;
  assign Accum2_acc_919_nl = nl_Accum2_acc_919_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1 = Accum2_acc_920_nl
      + Accum2_acc_919_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[949:945]));
  assign Product1_2_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1589:1585]));
  assign Product1_3_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_927_nl = (readslicef_20_16_4(Product1_2_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_927_nl = nl_Accum2_acc_927_nl[15:0];
  assign nl_Product1_4_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2229:2225]));
  assign Product1_4_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2869:2865]));
  assign Product1_5_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_926_nl = (readslicef_20_16_4(Product1_4_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_926_nl = nl_Accum2_acc_926_nl[15:0];
  assign nl_Product1_6_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3509:3505]));
  assign Product1_6_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4149:4145]));
  assign Product1_7_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_925_nl = (readslicef_20_16_4(Product1_6_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_925_nl = nl_Accum2_acc_925_nl[15:0];
  assign nl_Product1_8_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4789:4785]));
  assign Product1_8_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5429:5425]));
  assign Product1_9_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_924_nl = (readslicef_20_16_4(Product1_8_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_924_nl = nl_Accum2_acc_924_nl[15:0];
  assign nl_Accum2_acc_933_nl = Accum2_acc_927_nl + Accum2_acc_926_nl + Accum2_acc_925_nl
      + Accum2_acc_924_nl;
  assign Accum2_acc_933_nl = nl_Accum2_acc_933_nl[15:0];
  assign nl_Product1_10_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6069:6065]));
  assign Product1_10_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6709:6705]));
  assign Product1_11_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_923_nl = (readslicef_20_16_4(Product1_10_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_923_nl = nl_Accum2_acc_923_nl[15:0];
  assign nl_Product1_12_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7349:7345]));
  assign Product1_12_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7989:7985]));
  assign Product1_13_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_922_nl = (readslicef_20_16_4(Product1_12_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_922_nl = nl_Accum2_acc_922_nl[15:0];
  assign nl_Accum2_acc_929_nl = Accum2_acc_923_nl + Accum2_acc_922_nl;
  assign Accum2_acc_929_nl = nl_Accum2_acc_929_nl[15:0];
  assign nl_Accum2_acc_1853_nl = (Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[309:305]);
  assign Accum2_acc_1853_nl = nl_Accum2_acc_1853_nl[9:0];
  assign nl_Product1_1_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[309:305]));
  assign Product1_1_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_928_nl = ({Accum2_acc_1853_nl , (Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_928_nl = nl_Accum2_acc_928_nl[15:0];
  assign nl_Accum2_acc_932_nl = Accum2_acc_929_nl + Accum2_acc_928_nl;
  assign Accum2_acc_932_nl = nl_Accum2_acc_932_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1 = Accum2_acc_933_nl
      + Accum2_acc_932_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[954:950]));
  assign Product1_2_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1594:1590]));
  assign Product1_3_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_940_nl = (readslicef_20_16_4(Product1_2_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_940_nl = nl_Accum2_acc_940_nl[15:0];
  assign nl_Product1_4_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2234:2230]));
  assign Product1_4_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2874:2870]));
  assign Product1_5_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_939_nl = (readslicef_20_16_4(Product1_4_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_939_nl = nl_Accum2_acc_939_nl[15:0];
  assign nl_Product1_6_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3514:3510]));
  assign Product1_6_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4154:4150]));
  assign Product1_7_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_938_nl = (readslicef_20_16_4(Product1_6_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_938_nl = nl_Accum2_acc_938_nl[15:0];
  assign nl_Product1_8_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4794:4790]));
  assign Product1_8_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5434:5430]));
  assign Product1_9_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_937_nl = (readslicef_20_16_4(Product1_8_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_937_nl = nl_Accum2_acc_937_nl[15:0];
  assign nl_Accum2_acc_946_nl = Accum2_acc_940_nl + Accum2_acc_939_nl + Accum2_acc_938_nl
      + Accum2_acc_937_nl;
  assign Accum2_acc_946_nl = nl_Accum2_acc_946_nl[15:0];
  assign nl_Product1_10_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6074:6070]));
  assign Product1_10_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6714:6710]));
  assign Product1_11_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_936_nl = (readslicef_20_16_4(Product1_10_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_936_nl = nl_Accum2_acc_936_nl[15:0];
  assign nl_Product1_12_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7354:7350]));
  assign Product1_12_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7994:7990]));
  assign Product1_13_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_935_nl = (readslicef_20_16_4(Product1_12_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_935_nl = nl_Accum2_acc_935_nl[15:0];
  assign nl_Accum2_acc_942_nl = Accum2_acc_936_nl + Accum2_acc_935_nl;
  assign Accum2_acc_942_nl = nl_Accum2_acc_942_nl[15:0];
  assign nl_Accum2_acc_1854_nl = (Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[314:310]);
  assign Accum2_acc_1854_nl = nl_Accum2_acc_1854_nl[9:0];
  assign nl_Product1_1_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[314:310]));
  assign Product1_1_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_941_nl = ({Accum2_acc_1854_nl , (Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_941_nl = nl_Accum2_acc_941_nl[15:0];
  assign nl_Accum2_acc_945_nl = Accum2_acc_942_nl + Accum2_acc_941_nl;
  assign Accum2_acc_945_nl = nl_Accum2_acc_945_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1 = Accum2_acc_946_nl
      + Accum2_acc_945_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1 = (nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[959:955]));
  assign Product1_2_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1599:1595]));
  assign Product1_3_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_953_nl = (readslicef_20_16_4(Product1_2_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_953_nl = nl_Accum2_acc_953_nl[15:0];
  assign nl_Product1_4_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2239:2235]));
  assign Product1_4_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2879:2875]));
  assign Product1_5_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_952_nl = (readslicef_20_16_4(Product1_4_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_952_nl = nl_Accum2_acc_952_nl[15:0];
  assign nl_Product1_6_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3519:3515]));
  assign Product1_6_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4159:4155]));
  assign Product1_7_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_951_nl = (readslicef_20_16_4(Product1_6_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_951_nl = nl_Accum2_acc_951_nl[15:0];
  assign nl_Product1_8_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4799:4795]));
  assign Product1_8_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5439:5435]));
  assign Product1_9_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_950_nl = (readslicef_20_16_4(Product1_8_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_950_nl = nl_Accum2_acc_950_nl[15:0];
  assign nl_Accum2_acc_959_nl = Accum2_acc_953_nl + Accum2_acc_952_nl + Accum2_acc_951_nl
      + Accum2_acc_950_nl;
  assign Accum2_acc_959_nl = nl_Accum2_acc_959_nl[15:0];
  assign nl_Product1_10_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6079:6075]));
  assign Product1_10_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6719:6715]));
  assign Product1_11_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_949_nl = (readslicef_20_16_4(Product1_10_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_949_nl = nl_Accum2_acc_949_nl[15:0];
  assign nl_Product1_12_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7359:7355]));
  assign Product1_12_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[7999:7995]));
  assign Product1_13_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_948_nl = (readslicef_20_16_4(Product1_12_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_948_nl = nl_Accum2_acc_948_nl[15:0];
  assign nl_Accum2_acc_955_nl = Accum2_acc_949_nl + Accum2_acc_948_nl;
  assign Accum2_acc_955_nl = nl_Accum2_acc_955_nl[15:0];
  assign nl_Accum2_acc_1855_nl = (Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[319:315]);
  assign Accum2_acc_1855_nl = nl_Accum2_acc_1855_nl[9:0];
  assign nl_Product1_1_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[319:315]));
  assign Product1_1_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_954_nl = ({Accum2_acc_1855_nl , (Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_954_nl = nl_Accum2_acc_954_nl[15:0];
  assign nl_Accum2_acc_958_nl = Accum2_acc_955_nl + Accum2_acc_954_nl;
  assign Accum2_acc_958_nl = nl_Accum2_acc_958_nl[15:0];
  assign nl_nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1 = Accum2_acc_959_nl
      + Accum2_acc_958_nl;
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1 = nl_nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1 = (Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[964:960]));
  assign Product1_2_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1604:1600]));
  assign Product1_3_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_966_nl = (readslicef_20_16_4(Product1_2_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_966_nl = nl_Accum2_acc_966_nl[15:0];
  assign nl_Product1_4_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2244:2240]));
  assign Product1_4_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2884:2880]));
  assign Product1_5_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_965_nl = (readslicef_20_16_4(Product1_4_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_965_nl = nl_Accum2_acc_965_nl[15:0];
  assign nl_Product1_6_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3524:3520]));
  assign Product1_6_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4164:4160]));
  assign Product1_7_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_964_nl = (readslicef_20_16_4(Product1_6_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_964_nl = nl_Accum2_acc_964_nl[15:0];
  assign nl_Product1_8_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4804:4800]));
  assign Product1_8_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5444:5440]));
  assign Product1_9_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_963_nl = (readslicef_20_16_4(Product1_8_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_963_nl = nl_Accum2_acc_963_nl[15:0];
  assign nl_Accum2_acc_972_nl = Accum2_acc_966_nl + Accum2_acc_965_nl + Accum2_acc_964_nl
      + Accum2_acc_963_nl;
  assign Accum2_acc_972_nl = nl_Accum2_acc_972_nl[15:0];
  assign nl_Product1_10_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6084:6080]));
  assign Product1_10_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6724:6720]));
  assign Product1_11_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_962_nl = (readslicef_20_16_4(Product1_10_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_962_nl = nl_Accum2_acc_962_nl[15:0];
  assign nl_Product1_12_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7364:7360]));
  assign Product1_12_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8004:8000]));
  assign Product1_13_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_961_nl = (readslicef_20_16_4(Product1_12_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_961_nl = nl_Accum2_acc_961_nl[15:0];
  assign nl_Accum2_acc_968_nl = Accum2_acc_962_nl + Accum2_acc_961_nl;
  assign Accum2_acc_968_nl = nl_Accum2_acc_968_nl[15:0];
  assign nl_Accum2_acc_1856_nl = (Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[324:320]);
  assign Accum2_acc_1856_nl = nl_Accum2_acc_1856_nl[9:0];
  assign nl_Product1_1_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[324:320]));
  assign Product1_1_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_967_nl = ({Accum2_acc_1856_nl , (Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_967_nl = nl_Accum2_acc_967_nl[15:0];
  assign nl_Accum2_acc_971_nl = Accum2_acc_968_nl + Accum2_acc_967_nl;
  assign Accum2_acc_971_nl = nl_Accum2_acc_971_nl[15:0];
  assign nl_Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1 = Accum2_acc_972_nl + Accum2_acc_971_nl;
  assign Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1 = (Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[969:965]));
  assign Product1_2_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1609:1605]));
  assign Product1_3_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_979_nl = (readslicef_20_16_4(Product1_2_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_979_nl = nl_Accum2_acc_979_nl[15:0];
  assign nl_Product1_4_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2249:2245]));
  assign Product1_4_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2889:2885]));
  assign Product1_5_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_978_nl = (readslicef_20_16_4(Product1_4_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_978_nl = nl_Accum2_acc_978_nl[15:0];
  assign nl_Product1_6_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3529:3525]));
  assign Product1_6_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4169:4165]));
  assign Product1_7_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_977_nl = (readslicef_20_16_4(Product1_6_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_977_nl = nl_Accum2_acc_977_nl[15:0];
  assign nl_Product1_8_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4809:4805]));
  assign Product1_8_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5449:5445]));
  assign Product1_9_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_976_nl = (readslicef_20_16_4(Product1_8_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_976_nl = nl_Accum2_acc_976_nl[15:0];
  assign nl_Accum2_acc_985_nl = Accum2_acc_979_nl + Accum2_acc_978_nl + Accum2_acc_977_nl
      + Accum2_acc_976_nl;
  assign Accum2_acc_985_nl = nl_Accum2_acc_985_nl[15:0];
  assign nl_Product1_10_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6089:6085]));
  assign Product1_10_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6729:6725]));
  assign Product1_11_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_975_nl = (readslicef_20_16_4(Product1_10_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_975_nl = nl_Accum2_acc_975_nl[15:0];
  assign nl_Product1_12_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7369:7365]));
  assign Product1_12_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8009:8005]));
  assign Product1_13_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_974_nl = (readslicef_20_16_4(Product1_12_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_974_nl = nl_Accum2_acc_974_nl[15:0];
  assign nl_Accum2_acc_981_nl = Accum2_acc_975_nl + Accum2_acc_974_nl;
  assign Accum2_acc_981_nl = nl_Accum2_acc_981_nl[15:0];
  assign nl_Accum2_acc_1857_nl = (Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[329:325]);
  assign Accum2_acc_1857_nl = nl_Accum2_acc_1857_nl[9:0];
  assign nl_Product1_1_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[329:325]));
  assign Product1_1_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_980_nl = ({Accum2_acc_1857_nl , (Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_980_nl = nl_Accum2_acc_980_nl[15:0];
  assign nl_Accum2_acc_984_nl = Accum2_acc_981_nl + Accum2_acc_980_nl;
  assign Accum2_acc_984_nl = nl_Accum2_acc_984_nl[15:0];
  assign nl_Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1 = Accum2_acc_985_nl + Accum2_acc_984_nl;
  assign Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1 = (Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[974:970]));
  assign Product1_2_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1614:1610]));
  assign Product1_3_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_992_nl = (readslicef_20_16_4(Product1_2_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_992_nl = nl_Accum2_acc_992_nl[15:0];
  assign nl_Product1_4_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2254:2250]));
  assign Product1_4_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2894:2890]));
  assign Product1_5_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_991_nl = (readslicef_20_16_4(Product1_4_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_991_nl = nl_Accum2_acc_991_nl[15:0];
  assign nl_Product1_6_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3534:3530]));
  assign Product1_6_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4174:4170]));
  assign Product1_7_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_990_nl = (readslicef_20_16_4(Product1_6_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_990_nl = nl_Accum2_acc_990_nl[15:0];
  assign nl_Product1_8_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4814:4810]));
  assign Product1_8_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5454:5450]));
  assign Product1_9_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_989_nl = (readslicef_20_16_4(Product1_8_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_989_nl = nl_Accum2_acc_989_nl[15:0];
  assign nl_Accum2_acc_998_nl = Accum2_acc_992_nl + Accum2_acc_991_nl + Accum2_acc_990_nl
      + Accum2_acc_989_nl;
  assign Accum2_acc_998_nl = nl_Accum2_acc_998_nl[15:0];
  assign nl_Product1_10_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6094:6090]));
  assign Product1_10_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6734:6730]));
  assign Product1_11_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_988_nl = (readslicef_20_16_4(Product1_10_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_988_nl = nl_Accum2_acc_988_nl[15:0];
  assign nl_Product1_12_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7374:7370]));
  assign Product1_12_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8014:8010]));
  assign Product1_13_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_987_nl = (readslicef_20_16_4(Product1_12_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_987_nl = nl_Accum2_acc_987_nl[15:0];
  assign nl_Accum2_acc_994_nl = Accum2_acc_988_nl + Accum2_acc_987_nl;
  assign Accum2_acc_994_nl = nl_Accum2_acc_994_nl[15:0];
  assign nl_Accum2_acc_1858_nl = (Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[334:330]);
  assign Accum2_acc_1858_nl = nl_Accum2_acc_1858_nl[9:0];
  assign nl_Product1_1_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[334:330]));
  assign Product1_1_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_993_nl = ({Accum2_acc_1858_nl , (Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_993_nl = nl_Accum2_acc_993_nl[15:0];
  assign nl_Accum2_acc_997_nl = Accum2_acc_994_nl + Accum2_acc_993_nl;
  assign Accum2_acc_997_nl = nl_Accum2_acc_997_nl[15:0];
  assign nl_Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1 = Accum2_acc_998_nl + Accum2_acc_997_nl;
  assign Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1 = (Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[979:975]));
  assign Product1_2_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1619:1615]));
  assign Product1_3_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1005_nl = (readslicef_20_16_4(Product1_2_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1005_nl = nl_Accum2_acc_1005_nl[15:0];
  assign nl_Product1_4_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2259:2255]));
  assign Product1_4_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2899:2895]));
  assign Product1_5_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1004_nl = (readslicef_20_16_4(Product1_4_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1004_nl = nl_Accum2_acc_1004_nl[15:0];
  assign nl_Product1_6_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3539:3535]));
  assign Product1_6_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4179:4175]));
  assign Product1_7_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1003_nl = (readslicef_20_16_4(Product1_6_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1003_nl = nl_Accum2_acc_1003_nl[15:0];
  assign nl_Product1_8_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4819:4815]));
  assign Product1_8_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5459:5455]));
  assign Product1_9_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1002_nl = (readslicef_20_16_4(Product1_8_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1002_nl = nl_Accum2_acc_1002_nl[15:0];
  assign nl_Accum2_acc_1011_nl = Accum2_acc_1005_nl + Accum2_acc_1004_nl + Accum2_acc_1003_nl
      + Accum2_acc_1002_nl;
  assign Accum2_acc_1011_nl = nl_Accum2_acc_1011_nl[15:0];
  assign nl_Product1_10_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6099:6095]));
  assign Product1_10_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6739:6735]));
  assign Product1_11_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1001_nl = (readslicef_20_16_4(Product1_10_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1001_nl = nl_Accum2_acc_1001_nl[15:0];
  assign nl_Product1_12_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7379:7375]));
  assign Product1_12_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8019:8015]));
  assign Product1_13_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1000_nl = (readslicef_20_16_4(Product1_12_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1000_nl = nl_Accum2_acc_1000_nl[15:0];
  assign nl_Accum2_acc_1007_nl = Accum2_acc_1001_nl + Accum2_acc_1000_nl;
  assign Accum2_acc_1007_nl = nl_Accum2_acc_1007_nl[15:0];
  assign nl_Accum2_acc_1859_nl = (Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[339:335]);
  assign Accum2_acc_1859_nl = nl_Accum2_acc_1859_nl[9:0];
  assign nl_Product1_1_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[339:335]));
  assign Product1_1_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1006_nl = ({Accum2_acc_1859_nl , (Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1006_nl = nl_Accum2_acc_1006_nl[15:0];
  assign nl_Accum2_acc_1010_nl = Accum2_acc_1007_nl + Accum2_acc_1006_nl;
  assign Accum2_acc_1010_nl = nl_Accum2_acc_1010_nl[15:0];
  assign nl_Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1011_nl + Accum2_acc_1010_nl;
  assign Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1 = (Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[984:980]));
  assign Product1_2_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1624:1620]));
  assign Product1_3_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1018_nl = (readslicef_20_16_4(Product1_2_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1018_nl = nl_Accum2_acc_1018_nl[15:0];
  assign nl_Product1_4_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2264:2260]));
  assign Product1_4_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2904:2900]));
  assign Product1_5_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1017_nl = (readslicef_20_16_4(Product1_4_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1017_nl = nl_Accum2_acc_1017_nl[15:0];
  assign nl_Product1_6_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3544:3540]));
  assign Product1_6_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4184:4180]));
  assign Product1_7_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1016_nl = (readslicef_20_16_4(Product1_6_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1016_nl = nl_Accum2_acc_1016_nl[15:0];
  assign nl_Product1_8_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4824:4820]));
  assign Product1_8_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5464:5460]));
  assign Product1_9_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1015_nl = (readslicef_20_16_4(Product1_8_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1015_nl = nl_Accum2_acc_1015_nl[15:0];
  assign nl_Accum2_acc_1024_nl = Accum2_acc_1018_nl + Accum2_acc_1017_nl + Accum2_acc_1016_nl
      + Accum2_acc_1015_nl;
  assign Accum2_acc_1024_nl = nl_Accum2_acc_1024_nl[15:0];
  assign nl_Product1_10_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6104:6100]));
  assign Product1_10_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6744:6740]));
  assign Product1_11_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1014_nl = (readslicef_20_16_4(Product1_10_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1014_nl = nl_Accum2_acc_1014_nl[15:0];
  assign nl_Product1_12_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7384:7380]));
  assign Product1_12_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8024:8020]));
  assign Product1_13_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1013_nl = (readslicef_20_16_4(Product1_12_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1013_nl = nl_Accum2_acc_1013_nl[15:0];
  assign nl_Accum2_acc_1020_nl = Accum2_acc_1014_nl + Accum2_acc_1013_nl;
  assign Accum2_acc_1020_nl = nl_Accum2_acc_1020_nl[15:0];
  assign nl_Accum2_acc_1860_nl = (Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[344:340]);
  assign Accum2_acc_1860_nl = nl_Accum2_acc_1860_nl[9:0];
  assign nl_Product1_1_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[344:340]));
  assign Product1_1_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1019_nl = ({Accum2_acc_1860_nl , (Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1019_nl = nl_Accum2_acc_1019_nl[15:0];
  assign nl_Accum2_acc_1023_nl = Accum2_acc_1020_nl + Accum2_acc_1019_nl;
  assign Accum2_acc_1023_nl = nl_Accum2_acc_1023_nl[15:0];
  assign nl_Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1024_nl + Accum2_acc_1023_nl;
  assign Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1 = (Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[989:985]));
  assign Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1629:1625]));
  assign Product1_3_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1031_nl = (readslicef_20_16_4(Product1_2_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1031_nl = nl_Accum2_acc_1031_nl[15:0];
  assign nl_Product1_4_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2269:2265]));
  assign Product1_4_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2909:2905]));
  assign Product1_5_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1030_nl = (readslicef_20_16_4(Product1_4_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1030_nl = nl_Accum2_acc_1030_nl[15:0];
  assign nl_Product1_6_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3549:3545]));
  assign Product1_6_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4189:4185]));
  assign Product1_7_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1029_nl = (readslicef_20_16_4(Product1_6_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1029_nl = nl_Accum2_acc_1029_nl[15:0];
  assign nl_Product1_8_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4829:4825]));
  assign Product1_8_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5469:5465]));
  assign Product1_9_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1028_nl = (readslicef_20_16_4(Product1_8_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1028_nl = nl_Accum2_acc_1028_nl[15:0];
  assign nl_Accum2_acc_1037_nl = Accum2_acc_1031_nl + Accum2_acc_1030_nl + Accum2_acc_1029_nl
      + Accum2_acc_1028_nl;
  assign Accum2_acc_1037_nl = nl_Accum2_acc_1037_nl[15:0];
  assign nl_Product1_10_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6109:6105]));
  assign Product1_10_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6749:6745]));
  assign Product1_11_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1027_nl = (readslicef_20_16_4(Product1_10_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1027_nl = nl_Accum2_acc_1027_nl[15:0];
  assign nl_Product1_12_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7389:7385]));
  assign Product1_12_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8029:8025]));
  assign Product1_13_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1026_nl = (readslicef_20_16_4(Product1_12_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1026_nl = nl_Accum2_acc_1026_nl[15:0];
  assign nl_Accum2_acc_1033_nl = Accum2_acc_1027_nl + Accum2_acc_1026_nl;
  assign Accum2_acc_1033_nl = nl_Accum2_acc_1033_nl[15:0];
  assign nl_Accum2_acc_1861_nl = (Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[349:345]);
  assign Accum2_acc_1861_nl = nl_Accum2_acc_1861_nl[9:0];
  assign nl_Product1_1_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[349:345]));
  assign Product1_1_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1032_nl = ({Accum2_acc_1861_nl , (Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1032_nl = nl_Accum2_acc_1032_nl[15:0];
  assign nl_Accum2_acc_1036_nl = Accum2_acc_1033_nl + Accum2_acc_1032_nl;
  assign Accum2_acc_1036_nl = nl_Accum2_acc_1036_nl[15:0];
  assign nl_Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1037_nl + Accum2_acc_1036_nl;
  assign Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1 = (Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[994:990]));
  assign Product1_2_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1634:1630]));
  assign Product1_3_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1044_nl = (readslicef_20_16_4(Product1_2_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1044_nl = nl_Accum2_acc_1044_nl[15:0];
  assign nl_Product1_4_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2274:2270]));
  assign Product1_4_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2914:2910]));
  assign Product1_5_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1043_nl = (readslicef_20_16_4(Product1_4_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1043_nl = nl_Accum2_acc_1043_nl[15:0];
  assign nl_Product1_6_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3554:3550]));
  assign Product1_6_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4194:4190]));
  assign Product1_7_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1042_nl = (readslicef_20_16_4(Product1_6_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1042_nl = nl_Accum2_acc_1042_nl[15:0];
  assign nl_Product1_8_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4834:4830]));
  assign Product1_8_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5474:5470]));
  assign Product1_9_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1041_nl = (readslicef_20_16_4(Product1_8_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1041_nl = nl_Accum2_acc_1041_nl[15:0];
  assign nl_Accum2_acc_1050_nl = Accum2_acc_1044_nl + Accum2_acc_1043_nl + Accum2_acc_1042_nl
      + Accum2_acc_1041_nl;
  assign Accum2_acc_1050_nl = nl_Accum2_acc_1050_nl[15:0];
  assign nl_Product1_10_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6114:6110]));
  assign Product1_10_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6754:6750]));
  assign Product1_11_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1040_nl = (readslicef_20_16_4(Product1_10_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1040_nl = nl_Accum2_acc_1040_nl[15:0];
  assign nl_Product1_12_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7394:7390]));
  assign Product1_12_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8034:8030]));
  assign Product1_13_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1039_nl = (readslicef_20_16_4(Product1_12_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1039_nl = nl_Accum2_acc_1039_nl[15:0];
  assign nl_Accum2_acc_1046_nl = Accum2_acc_1040_nl + Accum2_acc_1039_nl;
  assign Accum2_acc_1046_nl = nl_Accum2_acc_1046_nl[15:0];
  assign nl_Accum2_acc_1862_nl = (Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[354:350]);
  assign Accum2_acc_1862_nl = nl_Accum2_acc_1862_nl[9:0];
  assign nl_Product1_1_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[354:350]));
  assign Product1_1_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1045_nl = ({Accum2_acc_1862_nl , (Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1045_nl = nl_Accum2_acc_1045_nl[15:0];
  assign nl_Accum2_acc_1049_nl = Accum2_acc_1046_nl + Accum2_acc_1045_nl;
  assign Accum2_acc_1049_nl = nl_Accum2_acc_1049_nl[15:0];
  assign nl_Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1050_nl + Accum2_acc_1049_nl;
  assign Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1 = (Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[999:995]));
  assign Product1_2_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1639:1635]));
  assign Product1_3_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1057_nl = (readslicef_20_16_4(Product1_2_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1057_nl = nl_Accum2_acc_1057_nl[15:0];
  assign nl_Product1_4_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2279:2275]));
  assign Product1_4_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2919:2915]));
  assign Product1_5_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1056_nl = (readslicef_20_16_4(Product1_4_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1056_nl = nl_Accum2_acc_1056_nl[15:0];
  assign nl_Product1_6_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3559:3555]));
  assign Product1_6_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4199:4195]));
  assign Product1_7_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1055_nl = (readslicef_20_16_4(Product1_6_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1055_nl = nl_Accum2_acc_1055_nl[15:0];
  assign nl_Product1_8_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4839:4835]));
  assign Product1_8_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5479:5475]));
  assign Product1_9_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1054_nl = (readslicef_20_16_4(Product1_8_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1054_nl = nl_Accum2_acc_1054_nl[15:0];
  assign nl_Accum2_acc_1063_nl = Accum2_acc_1057_nl + Accum2_acc_1056_nl + Accum2_acc_1055_nl
      + Accum2_acc_1054_nl;
  assign Accum2_acc_1063_nl = nl_Accum2_acc_1063_nl[15:0];
  assign nl_Product1_10_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6119:6115]));
  assign Product1_10_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6759:6755]));
  assign Product1_11_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1053_nl = (readslicef_20_16_4(Product1_10_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1053_nl = nl_Accum2_acc_1053_nl[15:0];
  assign nl_Product1_12_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7399:7395]));
  assign Product1_12_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8039:8035]));
  assign Product1_13_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1052_nl = (readslicef_20_16_4(Product1_12_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1052_nl = nl_Accum2_acc_1052_nl[15:0];
  assign nl_Accum2_acc_1059_nl = Accum2_acc_1053_nl + Accum2_acc_1052_nl;
  assign Accum2_acc_1059_nl = nl_Accum2_acc_1059_nl[15:0];
  assign nl_Accum2_acc_1863_nl = (Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[359:355]);
  assign Accum2_acc_1863_nl = nl_Accum2_acc_1863_nl[9:0];
  assign nl_Product1_1_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[359:355]));
  assign Product1_1_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1058_nl = ({Accum2_acc_1863_nl , (Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1058_nl = nl_Accum2_acc_1058_nl[15:0];
  assign nl_Accum2_acc_1062_nl = Accum2_acc_1059_nl + Accum2_acc_1058_nl;
  assign Accum2_acc_1062_nl = nl_Accum2_acc_1062_nl[15:0];
  assign nl_Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1063_nl + Accum2_acc_1062_nl;
  assign Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1 = (Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1004:1000]));
  assign Product1_2_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1644:1640]));
  assign Product1_3_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1070_nl = (readslicef_20_16_4(Product1_2_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1070_nl = nl_Accum2_acc_1070_nl[15:0];
  assign nl_Product1_4_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2284:2280]));
  assign Product1_4_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2924:2920]));
  assign Product1_5_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1069_nl = (readslicef_20_16_4(Product1_4_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1069_nl = nl_Accum2_acc_1069_nl[15:0];
  assign nl_Product1_6_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3564:3560]));
  assign Product1_6_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4204:4200]));
  assign Product1_7_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1068_nl = (readslicef_20_16_4(Product1_6_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1068_nl = nl_Accum2_acc_1068_nl[15:0];
  assign nl_Product1_8_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4844:4840]));
  assign Product1_8_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5484:5480]));
  assign Product1_9_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1067_nl = (readslicef_20_16_4(Product1_8_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1067_nl = nl_Accum2_acc_1067_nl[15:0];
  assign nl_Accum2_acc_1076_nl = Accum2_acc_1070_nl + Accum2_acc_1069_nl + Accum2_acc_1068_nl
      + Accum2_acc_1067_nl;
  assign Accum2_acc_1076_nl = nl_Accum2_acc_1076_nl[15:0];
  assign nl_Product1_10_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6124:6120]));
  assign Product1_10_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6764:6760]));
  assign Product1_11_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1066_nl = (readslicef_20_16_4(Product1_10_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1066_nl = nl_Accum2_acc_1066_nl[15:0];
  assign nl_Product1_12_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7404:7400]));
  assign Product1_12_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8044:8040]));
  assign Product1_13_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1065_nl = (readslicef_20_16_4(Product1_12_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1065_nl = nl_Accum2_acc_1065_nl[15:0];
  assign nl_Accum2_acc_1072_nl = Accum2_acc_1066_nl + Accum2_acc_1065_nl;
  assign Accum2_acc_1072_nl = nl_Accum2_acc_1072_nl[15:0];
  assign nl_Accum2_acc_1864_nl = (Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[364:360]);
  assign Accum2_acc_1864_nl = nl_Accum2_acc_1864_nl[9:0];
  assign nl_Product1_1_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[364:360]));
  assign Product1_1_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1071_nl = ({Accum2_acc_1864_nl , (Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1071_nl = nl_Accum2_acc_1071_nl[15:0];
  assign nl_Accum2_acc_1075_nl = Accum2_acc_1072_nl + Accum2_acc_1071_nl;
  assign Accum2_acc_1075_nl = nl_Accum2_acc_1075_nl[15:0];
  assign nl_Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1076_nl + Accum2_acc_1075_nl;
  assign Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1 = (Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1009:1005]));
  assign Product1_2_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1649:1645]));
  assign Product1_3_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1083_nl = (readslicef_20_16_4(Product1_2_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1083_nl = nl_Accum2_acc_1083_nl[15:0];
  assign nl_Product1_4_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2289:2285]));
  assign Product1_4_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2929:2925]));
  assign Product1_5_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1082_nl = (readslicef_20_16_4(Product1_4_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1082_nl = nl_Accum2_acc_1082_nl[15:0];
  assign nl_Product1_6_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3569:3565]));
  assign Product1_6_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4209:4205]));
  assign Product1_7_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1081_nl = (readslicef_20_16_4(Product1_6_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1081_nl = nl_Accum2_acc_1081_nl[15:0];
  assign nl_Product1_8_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4849:4845]));
  assign Product1_8_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5489:5485]));
  assign Product1_9_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1080_nl = (readslicef_20_16_4(Product1_8_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1080_nl = nl_Accum2_acc_1080_nl[15:0];
  assign nl_Accum2_acc_1089_nl = Accum2_acc_1083_nl + Accum2_acc_1082_nl + Accum2_acc_1081_nl
      + Accum2_acc_1080_nl;
  assign Accum2_acc_1089_nl = nl_Accum2_acc_1089_nl[15:0];
  assign nl_Product1_10_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6129:6125]));
  assign Product1_10_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6769:6765]));
  assign Product1_11_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1079_nl = (readslicef_20_16_4(Product1_10_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1079_nl = nl_Accum2_acc_1079_nl[15:0];
  assign nl_Product1_12_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7409:7405]));
  assign Product1_12_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8049:8045]));
  assign Product1_13_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1078_nl = (readslicef_20_16_4(Product1_12_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1078_nl = nl_Accum2_acc_1078_nl[15:0];
  assign nl_Accum2_acc_1085_nl = Accum2_acc_1079_nl + Accum2_acc_1078_nl;
  assign Accum2_acc_1085_nl = nl_Accum2_acc_1085_nl[15:0];
  assign nl_Accum2_acc_1865_nl = (Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[369:365]);
  assign Accum2_acc_1865_nl = nl_Accum2_acc_1865_nl[9:0];
  assign nl_Product1_1_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[369:365]));
  assign Product1_1_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1084_nl = ({Accum2_acc_1865_nl , (Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1084_nl = nl_Accum2_acc_1084_nl[15:0];
  assign nl_Accum2_acc_1088_nl = Accum2_acc_1085_nl + Accum2_acc_1084_nl;
  assign Accum2_acc_1088_nl = nl_Accum2_acc_1088_nl[15:0];
  assign nl_Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1089_nl + Accum2_acc_1088_nl;
  assign Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1 = (Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1014:1010]));
  assign Product1_2_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1654:1650]));
  assign Product1_3_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1096_nl = (readslicef_20_16_4(Product1_2_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1096_nl = nl_Accum2_acc_1096_nl[15:0];
  assign nl_Product1_4_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2294:2290]));
  assign Product1_4_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2934:2930]));
  assign Product1_5_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1095_nl = (readslicef_20_16_4(Product1_4_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1095_nl = nl_Accum2_acc_1095_nl[15:0];
  assign nl_Product1_6_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3574:3570]));
  assign Product1_6_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4214:4210]));
  assign Product1_7_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1094_nl = (readslicef_20_16_4(Product1_6_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1094_nl = nl_Accum2_acc_1094_nl[15:0];
  assign nl_Product1_8_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4854:4850]));
  assign Product1_8_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5494:5490]));
  assign Product1_9_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1093_nl = (readslicef_20_16_4(Product1_8_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1093_nl = nl_Accum2_acc_1093_nl[15:0];
  assign nl_Accum2_acc_1102_nl = Accum2_acc_1096_nl + Accum2_acc_1095_nl + Accum2_acc_1094_nl
      + Accum2_acc_1093_nl;
  assign Accum2_acc_1102_nl = nl_Accum2_acc_1102_nl[15:0];
  assign nl_Product1_10_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6134:6130]));
  assign Product1_10_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6774:6770]));
  assign Product1_11_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1092_nl = (readslicef_20_16_4(Product1_10_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1092_nl = nl_Accum2_acc_1092_nl[15:0];
  assign nl_Product1_12_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7414:7410]));
  assign Product1_12_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8054:8050]));
  assign Product1_13_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1091_nl = (readslicef_20_16_4(Product1_12_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1091_nl = nl_Accum2_acc_1091_nl[15:0];
  assign nl_Accum2_acc_1098_nl = Accum2_acc_1092_nl + Accum2_acc_1091_nl;
  assign Accum2_acc_1098_nl = nl_Accum2_acc_1098_nl[15:0];
  assign nl_Accum2_acc_1866_nl = (Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[374:370]);
  assign Accum2_acc_1866_nl = nl_Accum2_acc_1866_nl[9:0];
  assign nl_Product1_1_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[374:370]));
  assign Product1_1_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1097_nl = ({Accum2_acc_1866_nl , (Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1097_nl = nl_Accum2_acc_1097_nl[15:0];
  assign nl_Accum2_acc_1101_nl = Accum2_acc_1098_nl + Accum2_acc_1097_nl;
  assign Accum2_acc_1101_nl = nl_Accum2_acc_1101_nl[15:0];
  assign nl_Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1102_nl + Accum2_acc_1101_nl;
  assign Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1 = (Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1019:1015]));
  assign Product1_2_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1659:1655]));
  assign Product1_3_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1109_nl = (readslicef_20_16_4(Product1_2_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1109_nl = nl_Accum2_acc_1109_nl[15:0];
  assign nl_Product1_4_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2299:2295]));
  assign Product1_4_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2939:2935]));
  assign Product1_5_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1108_nl = (readslicef_20_16_4(Product1_4_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1108_nl = nl_Accum2_acc_1108_nl[15:0];
  assign nl_Product1_6_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3579:3575]));
  assign Product1_6_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4219:4215]));
  assign Product1_7_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1107_nl = (readslicef_20_16_4(Product1_6_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1107_nl = nl_Accum2_acc_1107_nl[15:0];
  assign nl_Product1_8_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4859:4855]));
  assign Product1_8_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5499:5495]));
  assign Product1_9_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1106_nl = (readslicef_20_16_4(Product1_8_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1106_nl = nl_Accum2_acc_1106_nl[15:0];
  assign nl_Accum2_acc_1115_nl = Accum2_acc_1109_nl + Accum2_acc_1108_nl + Accum2_acc_1107_nl
      + Accum2_acc_1106_nl;
  assign Accum2_acc_1115_nl = nl_Accum2_acc_1115_nl[15:0];
  assign nl_Product1_10_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6139:6135]));
  assign Product1_10_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6779:6775]));
  assign Product1_11_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1105_nl = (readslicef_20_16_4(Product1_10_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1105_nl = nl_Accum2_acc_1105_nl[15:0];
  assign nl_Product1_12_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7419:7415]));
  assign Product1_12_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8059:8055]));
  assign Product1_13_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1104_nl = (readslicef_20_16_4(Product1_12_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1104_nl = nl_Accum2_acc_1104_nl[15:0];
  assign nl_Accum2_acc_1111_nl = Accum2_acc_1105_nl + Accum2_acc_1104_nl;
  assign Accum2_acc_1111_nl = nl_Accum2_acc_1111_nl[15:0];
  assign nl_Accum2_acc_1867_nl = (Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[379:375]);
  assign Accum2_acc_1867_nl = nl_Accum2_acc_1867_nl[9:0];
  assign nl_Product1_1_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[379:375]));
  assign Product1_1_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1110_nl = ({Accum2_acc_1867_nl , (Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1110_nl = nl_Accum2_acc_1110_nl[15:0];
  assign nl_Accum2_acc_1114_nl = Accum2_acc_1111_nl + Accum2_acc_1110_nl;
  assign Accum2_acc_1114_nl = nl_Accum2_acc_1114_nl[15:0];
  assign nl_Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1115_nl + Accum2_acc_1114_nl;
  assign Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1 = (Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1024:1020]));
  assign Product1_2_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1664:1660]));
  assign Product1_3_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1122_nl = (readslicef_20_16_4(Product1_2_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1122_nl = nl_Accum2_acc_1122_nl[15:0];
  assign nl_Product1_4_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2304:2300]));
  assign Product1_4_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2944:2940]));
  assign Product1_5_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1121_nl = (readslicef_20_16_4(Product1_4_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1121_nl = nl_Accum2_acc_1121_nl[15:0];
  assign nl_Product1_6_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3584:3580]));
  assign Product1_6_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4224:4220]));
  assign Product1_7_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1120_nl = (readslicef_20_16_4(Product1_6_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1120_nl = nl_Accum2_acc_1120_nl[15:0];
  assign nl_Product1_8_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4864:4860]));
  assign Product1_8_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5504:5500]));
  assign Product1_9_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1119_nl = (readslicef_20_16_4(Product1_8_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1119_nl = nl_Accum2_acc_1119_nl[15:0];
  assign nl_Accum2_acc_1128_nl = Accum2_acc_1122_nl + Accum2_acc_1121_nl + Accum2_acc_1120_nl
      + Accum2_acc_1119_nl;
  assign Accum2_acc_1128_nl = nl_Accum2_acc_1128_nl[15:0];
  assign nl_Product1_10_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6144:6140]));
  assign Product1_10_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6784:6780]));
  assign Product1_11_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1118_nl = (readslicef_20_16_4(Product1_10_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1118_nl = nl_Accum2_acc_1118_nl[15:0];
  assign nl_Product1_12_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7424:7420]));
  assign Product1_12_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8064:8060]));
  assign Product1_13_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1117_nl = (readslicef_20_16_4(Product1_12_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1117_nl = nl_Accum2_acc_1117_nl[15:0];
  assign nl_Accum2_acc_1124_nl = Accum2_acc_1118_nl + Accum2_acc_1117_nl;
  assign Accum2_acc_1124_nl = nl_Accum2_acc_1124_nl[15:0];
  assign nl_Accum2_acc_1868_nl = (Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[384:380]);
  assign Accum2_acc_1868_nl = nl_Accum2_acc_1868_nl[9:0];
  assign nl_Product1_1_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[384:380]));
  assign Product1_1_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1123_nl = ({Accum2_acc_1868_nl , (Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1123_nl = nl_Accum2_acc_1123_nl[15:0];
  assign nl_Accum2_acc_1127_nl = Accum2_acc_1124_nl + Accum2_acc_1123_nl;
  assign Accum2_acc_1127_nl = nl_Accum2_acc_1127_nl[15:0];
  assign nl_Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1128_nl + Accum2_acc_1127_nl;
  assign Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1 = (Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1029:1025]));
  assign Product1_2_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1669:1665]));
  assign Product1_3_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1135_nl = (readslicef_20_16_4(Product1_2_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1135_nl = nl_Accum2_acc_1135_nl[15:0];
  assign nl_Product1_4_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2309:2305]));
  assign Product1_4_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2949:2945]));
  assign Product1_5_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1134_nl = (readslicef_20_16_4(Product1_4_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1134_nl = nl_Accum2_acc_1134_nl[15:0];
  assign nl_Product1_6_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3589:3585]));
  assign Product1_6_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4229:4225]));
  assign Product1_7_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1133_nl = (readslicef_20_16_4(Product1_6_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1133_nl = nl_Accum2_acc_1133_nl[15:0];
  assign nl_Product1_8_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4869:4865]));
  assign Product1_8_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5509:5505]));
  assign Product1_9_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1132_nl = (readslicef_20_16_4(Product1_8_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1132_nl = nl_Accum2_acc_1132_nl[15:0];
  assign nl_Accum2_acc_1141_nl = Accum2_acc_1135_nl + Accum2_acc_1134_nl + Accum2_acc_1133_nl
      + Accum2_acc_1132_nl;
  assign Accum2_acc_1141_nl = nl_Accum2_acc_1141_nl[15:0];
  assign nl_Product1_10_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6149:6145]));
  assign Product1_10_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6789:6785]));
  assign Product1_11_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1131_nl = (readslicef_20_16_4(Product1_10_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1131_nl = nl_Accum2_acc_1131_nl[15:0];
  assign nl_Product1_12_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7429:7425]));
  assign Product1_12_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8069:8065]));
  assign Product1_13_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1130_nl = (readslicef_20_16_4(Product1_12_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1130_nl = nl_Accum2_acc_1130_nl[15:0];
  assign nl_Accum2_acc_1137_nl = Accum2_acc_1131_nl + Accum2_acc_1130_nl;
  assign Accum2_acc_1137_nl = nl_Accum2_acc_1137_nl[15:0];
  assign nl_Accum2_acc_1869_nl = (Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[389:385]);
  assign Accum2_acc_1869_nl = nl_Accum2_acc_1869_nl[9:0];
  assign nl_Product1_1_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[389:385]));
  assign Product1_1_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1136_nl = ({Accum2_acc_1869_nl , (Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1136_nl = nl_Accum2_acc_1136_nl[15:0];
  assign nl_Accum2_acc_1140_nl = Accum2_acc_1137_nl + Accum2_acc_1136_nl;
  assign Accum2_acc_1140_nl = nl_Accum2_acc_1140_nl[15:0];
  assign nl_Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1141_nl + Accum2_acc_1140_nl;
  assign Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1 = (Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1034:1030]));
  assign Product1_2_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1674:1670]));
  assign Product1_3_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1148_nl = (readslicef_20_16_4(Product1_2_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1148_nl = nl_Accum2_acc_1148_nl[15:0];
  assign nl_Product1_4_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2314:2310]));
  assign Product1_4_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2954:2950]));
  assign Product1_5_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1147_nl = (readslicef_20_16_4(Product1_4_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1147_nl = nl_Accum2_acc_1147_nl[15:0];
  assign nl_Product1_6_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3594:3590]));
  assign Product1_6_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4234:4230]));
  assign Product1_7_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1146_nl = (readslicef_20_16_4(Product1_6_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1146_nl = nl_Accum2_acc_1146_nl[15:0];
  assign nl_Product1_8_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4874:4870]));
  assign Product1_8_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5514:5510]));
  assign Product1_9_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1145_nl = (readslicef_20_16_4(Product1_8_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1145_nl = nl_Accum2_acc_1145_nl[15:0];
  assign nl_Accum2_acc_1154_nl = Accum2_acc_1148_nl + Accum2_acc_1147_nl + Accum2_acc_1146_nl
      + Accum2_acc_1145_nl;
  assign Accum2_acc_1154_nl = nl_Accum2_acc_1154_nl[15:0];
  assign nl_Product1_10_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6154:6150]));
  assign Product1_10_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6794:6790]));
  assign Product1_11_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1144_nl = (readslicef_20_16_4(Product1_10_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1144_nl = nl_Accum2_acc_1144_nl[15:0];
  assign nl_Product1_12_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7434:7430]));
  assign Product1_12_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8074:8070]));
  assign Product1_13_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1143_nl = (readslicef_20_16_4(Product1_12_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1143_nl = nl_Accum2_acc_1143_nl[15:0];
  assign nl_Accum2_acc_1150_nl = Accum2_acc_1144_nl + Accum2_acc_1143_nl;
  assign Accum2_acc_1150_nl = nl_Accum2_acc_1150_nl[15:0];
  assign nl_Accum2_acc_1870_nl = (Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[394:390]);
  assign Accum2_acc_1870_nl = nl_Accum2_acc_1870_nl[9:0];
  assign nl_Product1_1_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[394:390]));
  assign Product1_1_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1149_nl = ({Accum2_acc_1870_nl , (Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1149_nl = nl_Accum2_acc_1149_nl[15:0];
  assign nl_Accum2_acc_1153_nl = Accum2_acc_1150_nl + Accum2_acc_1149_nl;
  assign Accum2_acc_1153_nl = nl_Accum2_acc_1153_nl[15:0];
  assign nl_Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1154_nl + Accum2_acc_1153_nl;
  assign Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1 = (Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1039:1035]));
  assign Product1_2_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1679:1675]));
  assign Product1_3_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1161_nl = (readslicef_20_16_4(Product1_2_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1161_nl = nl_Accum2_acc_1161_nl[15:0];
  assign nl_Product1_4_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2319:2315]));
  assign Product1_4_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2959:2955]));
  assign Product1_5_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1160_nl = (readslicef_20_16_4(Product1_4_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1160_nl = nl_Accum2_acc_1160_nl[15:0];
  assign nl_Product1_6_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3599:3595]));
  assign Product1_6_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4239:4235]));
  assign Product1_7_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1159_nl = (readslicef_20_16_4(Product1_6_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1159_nl = nl_Accum2_acc_1159_nl[15:0];
  assign nl_Product1_8_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4879:4875]));
  assign Product1_8_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5519:5515]));
  assign Product1_9_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1158_nl = (readslicef_20_16_4(Product1_8_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1158_nl = nl_Accum2_acc_1158_nl[15:0];
  assign nl_Accum2_acc_1167_nl = Accum2_acc_1161_nl + Accum2_acc_1160_nl + Accum2_acc_1159_nl
      + Accum2_acc_1158_nl;
  assign Accum2_acc_1167_nl = nl_Accum2_acc_1167_nl[15:0];
  assign nl_Product1_10_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6159:6155]));
  assign Product1_10_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6799:6795]));
  assign Product1_11_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1157_nl = (readslicef_20_16_4(Product1_10_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1157_nl = nl_Accum2_acc_1157_nl[15:0];
  assign nl_Product1_12_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7439:7435]));
  assign Product1_12_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8079:8075]));
  assign Product1_13_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1156_nl = (readslicef_20_16_4(Product1_12_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1156_nl = nl_Accum2_acc_1156_nl[15:0];
  assign nl_Accum2_acc_1163_nl = Accum2_acc_1157_nl + Accum2_acc_1156_nl;
  assign Accum2_acc_1163_nl = nl_Accum2_acc_1163_nl[15:0];
  assign nl_Accum2_acc_1871_nl = (Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[399:395]);
  assign Accum2_acc_1871_nl = nl_Accum2_acc_1871_nl[9:0];
  assign nl_Product1_1_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[399:395]));
  assign Product1_1_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1162_nl = ({Accum2_acc_1871_nl , (Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1162_nl = nl_Accum2_acc_1162_nl[15:0];
  assign nl_Accum2_acc_1166_nl = Accum2_acc_1163_nl + Accum2_acc_1162_nl;
  assign Accum2_acc_1166_nl = nl_Accum2_acc_1166_nl[15:0];
  assign nl_Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1167_nl + Accum2_acc_1166_nl;
  assign Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1 = (Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1044:1040]));
  assign Product1_2_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1684:1680]));
  assign Product1_3_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1174_nl = (readslicef_20_16_4(Product1_2_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1174_nl = nl_Accum2_acc_1174_nl[15:0];
  assign nl_Product1_4_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2324:2320]));
  assign Product1_4_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2964:2960]));
  assign Product1_5_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1173_nl = (readslicef_20_16_4(Product1_4_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1173_nl = nl_Accum2_acc_1173_nl[15:0];
  assign nl_Product1_6_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3604:3600]));
  assign Product1_6_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4244:4240]));
  assign Product1_7_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1172_nl = (readslicef_20_16_4(Product1_6_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1172_nl = nl_Accum2_acc_1172_nl[15:0];
  assign nl_Product1_8_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4884:4880]));
  assign Product1_8_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5524:5520]));
  assign Product1_9_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1171_nl = (readslicef_20_16_4(Product1_8_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1171_nl = nl_Accum2_acc_1171_nl[15:0];
  assign nl_Accum2_acc_1180_nl = Accum2_acc_1174_nl + Accum2_acc_1173_nl + Accum2_acc_1172_nl
      + Accum2_acc_1171_nl;
  assign Accum2_acc_1180_nl = nl_Accum2_acc_1180_nl[15:0];
  assign nl_Product1_10_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6164:6160]));
  assign Product1_10_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6804:6800]));
  assign Product1_11_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1170_nl = (readslicef_20_16_4(Product1_10_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1170_nl = nl_Accum2_acc_1170_nl[15:0];
  assign nl_Product1_12_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7444:7440]));
  assign Product1_12_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8084:8080]));
  assign Product1_13_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1169_nl = (readslicef_20_16_4(Product1_12_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1169_nl = nl_Accum2_acc_1169_nl[15:0];
  assign nl_Accum2_acc_1176_nl = Accum2_acc_1170_nl + Accum2_acc_1169_nl;
  assign Accum2_acc_1176_nl = nl_Accum2_acc_1176_nl[15:0];
  assign nl_Accum2_acc_1872_nl = (Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[404:400]);
  assign Accum2_acc_1872_nl = nl_Accum2_acc_1872_nl[9:0];
  assign nl_Product1_1_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[404:400]));
  assign Product1_1_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1175_nl = ({Accum2_acc_1872_nl , (Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1175_nl = nl_Accum2_acc_1175_nl[15:0];
  assign nl_Accum2_acc_1179_nl = Accum2_acc_1176_nl + Accum2_acc_1175_nl;
  assign Accum2_acc_1179_nl = nl_Accum2_acc_1179_nl[15:0];
  assign nl_Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1180_nl + Accum2_acc_1179_nl;
  assign Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1 = (Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1049:1045]));
  assign Product1_2_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1689:1685]));
  assign Product1_3_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1187_nl = (readslicef_20_16_4(Product1_2_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1187_nl = nl_Accum2_acc_1187_nl[15:0];
  assign nl_Product1_4_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2329:2325]));
  assign Product1_4_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2969:2965]));
  assign Product1_5_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1186_nl = (readslicef_20_16_4(Product1_4_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1186_nl = nl_Accum2_acc_1186_nl[15:0];
  assign nl_Product1_6_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3609:3605]));
  assign Product1_6_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4249:4245]));
  assign Product1_7_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1185_nl = (readslicef_20_16_4(Product1_6_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1185_nl = nl_Accum2_acc_1185_nl[15:0];
  assign nl_Product1_8_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4889:4885]));
  assign Product1_8_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5529:5525]));
  assign Product1_9_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1184_nl = (readslicef_20_16_4(Product1_8_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1184_nl = nl_Accum2_acc_1184_nl[15:0];
  assign nl_Accum2_acc_1193_nl = Accum2_acc_1187_nl + Accum2_acc_1186_nl + Accum2_acc_1185_nl
      + Accum2_acc_1184_nl;
  assign Accum2_acc_1193_nl = nl_Accum2_acc_1193_nl[15:0];
  assign nl_Product1_10_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6169:6165]));
  assign Product1_10_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6809:6805]));
  assign Product1_11_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1183_nl = (readslicef_20_16_4(Product1_10_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1183_nl = nl_Accum2_acc_1183_nl[15:0];
  assign nl_Product1_12_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7449:7445]));
  assign Product1_12_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8089:8085]));
  assign Product1_13_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1182_nl = (readslicef_20_16_4(Product1_12_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1182_nl = nl_Accum2_acc_1182_nl[15:0];
  assign nl_Accum2_acc_1189_nl = Accum2_acc_1183_nl + Accum2_acc_1182_nl;
  assign Accum2_acc_1189_nl = nl_Accum2_acc_1189_nl[15:0];
  assign nl_Accum2_acc_1873_nl = (Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[409:405]);
  assign Accum2_acc_1873_nl = nl_Accum2_acc_1873_nl[9:0];
  assign nl_Product1_1_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[409:405]));
  assign Product1_1_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1188_nl = ({Accum2_acc_1873_nl , (Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1188_nl = nl_Accum2_acc_1188_nl[15:0];
  assign nl_Accum2_acc_1192_nl = Accum2_acc_1189_nl + Accum2_acc_1188_nl;
  assign Accum2_acc_1192_nl = nl_Accum2_acc_1192_nl[15:0];
  assign nl_Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1193_nl + Accum2_acc_1192_nl;
  assign Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1 = (Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1054:1050]));
  assign Product1_2_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1694:1690]));
  assign Product1_3_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1200_nl = (readslicef_20_16_4(Product1_2_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1200_nl = nl_Accum2_acc_1200_nl[15:0];
  assign nl_Product1_4_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2334:2330]));
  assign Product1_4_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2974:2970]));
  assign Product1_5_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1199_nl = (readslicef_20_16_4(Product1_4_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1199_nl = nl_Accum2_acc_1199_nl[15:0];
  assign nl_Product1_6_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3614:3610]));
  assign Product1_6_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4254:4250]));
  assign Product1_7_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1198_nl = (readslicef_20_16_4(Product1_6_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1198_nl = nl_Accum2_acc_1198_nl[15:0];
  assign nl_Product1_8_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4894:4890]));
  assign Product1_8_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5534:5530]));
  assign Product1_9_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1197_nl = (readslicef_20_16_4(Product1_8_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1197_nl = nl_Accum2_acc_1197_nl[15:0];
  assign nl_Accum2_acc_1206_nl = Accum2_acc_1200_nl + Accum2_acc_1199_nl + Accum2_acc_1198_nl
      + Accum2_acc_1197_nl;
  assign Accum2_acc_1206_nl = nl_Accum2_acc_1206_nl[15:0];
  assign nl_Product1_10_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6174:6170]));
  assign Product1_10_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6814:6810]));
  assign Product1_11_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1196_nl = (readslicef_20_16_4(Product1_10_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1196_nl = nl_Accum2_acc_1196_nl[15:0];
  assign nl_Product1_12_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7454:7450]));
  assign Product1_12_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8094:8090]));
  assign Product1_13_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1195_nl = (readslicef_20_16_4(Product1_12_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1195_nl = nl_Accum2_acc_1195_nl[15:0];
  assign nl_Accum2_acc_1202_nl = Accum2_acc_1196_nl + Accum2_acc_1195_nl;
  assign Accum2_acc_1202_nl = nl_Accum2_acc_1202_nl[15:0];
  assign nl_Accum2_acc_1874_nl = (Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[414:410]);
  assign Accum2_acc_1874_nl = nl_Accum2_acc_1874_nl[9:0];
  assign nl_Product1_1_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[414:410]));
  assign Product1_1_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1201_nl = ({Accum2_acc_1874_nl , (Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1201_nl = nl_Accum2_acc_1201_nl[15:0];
  assign nl_Accum2_acc_1205_nl = Accum2_acc_1202_nl + Accum2_acc_1201_nl;
  assign Accum2_acc_1205_nl = nl_Accum2_acc_1205_nl[15:0];
  assign nl_Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1206_nl + Accum2_acc_1205_nl;
  assign Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1 = (Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1059:1055]));
  assign Product1_2_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1699:1695]));
  assign Product1_3_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1213_nl = (readslicef_20_16_4(Product1_2_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1213_nl = nl_Accum2_acc_1213_nl[15:0];
  assign nl_Product1_4_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2339:2335]));
  assign Product1_4_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2979:2975]));
  assign Product1_5_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1212_nl = (readslicef_20_16_4(Product1_4_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1212_nl = nl_Accum2_acc_1212_nl[15:0];
  assign nl_Product1_6_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3619:3615]));
  assign Product1_6_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4259:4255]));
  assign Product1_7_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1211_nl = (readslicef_20_16_4(Product1_6_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1211_nl = nl_Accum2_acc_1211_nl[15:0];
  assign nl_Product1_8_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4899:4895]));
  assign Product1_8_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5539:5535]));
  assign Product1_9_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1210_nl = (readslicef_20_16_4(Product1_8_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1210_nl = nl_Accum2_acc_1210_nl[15:0];
  assign nl_Accum2_acc_1219_nl = Accum2_acc_1213_nl + Accum2_acc_1212_nl + Accum2_acc_1211_nl
      + Accum2_acc_1210_nl;
  assign Accum2_acc_1219_nl = nl_Accum2_acc_1219_nl[15:0];
  assign nl_Product1_10_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6179:6175]));
  assign Product1_10_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6819:6815]));
  assign Product1_11_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1209_nl = (readslicef_20_16_4(Product1_10_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1209_nl = nl_Accum2_acc_1209_nl[15:0];
  assign nl_Product1_12_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7459:7455]));
  assign Product1_12_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8099:8095]));
  assign Product1_13_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1208_nl = (readslicef_20_16_4(Product1_12_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1208_nl = nl_Accum2_acc_1208_nl[15:0];
  assign nl_Accum2_acc_1215_nl = Accum2_acc_1209_nl + Accum2_acc_1208_nl;
  assign Accum2_acc_1215_nl = nl_Accum2_acc_1215_nl[15:0];
  assign nl_Accum2_acc_1875_nl = (Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[419:415]);
  assign Accum2_acc_1875_nl = nl_Accum2_acc_1875_nl[9:0];
  assign nl_Product1_1_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[419:415]));
  assign Product1_1_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1214_nl = ({Accum2_acc_1875_nl , (Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1214_nl = nl_Accum2_acc_1214_nl[15:0];
  assign nl_Accum2_acc_1218_nl = Accum2_acc_1215_nl + Accum2_acc_1214_nl;
  assign Accum2_acc_1218_nl = nl_Accum2_acc_1218_nl[15:0];
  assign nl_Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1219_nl + Accum2_acc_1218_nl;
  assign Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1 = (Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1064:1060]));
  assign Product1_2_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1704:1700]));
  assign Product1_3_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1226_nl = (readslicef_20_16_4(Product1_2_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1226_nl = nl_Accum2_acc_1226_nl[15:0];
  assign nl_Product1_4_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2344:2340]));
  assign Product1_4_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2984:2980]));
  assign Product1_5_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1225_nl = (readslicef_20_16_4(Product1_4_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1225_nl = nl_Accum2_acc_1225_nl[15:0];
  assign nl_Product1_6_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3624:3620]));
  assign Product1_6_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4264:4260]));
  assign Product1_7_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1224_nl = (readslicef_20_16_4(Product1_6_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1224_nl = nl_Accum2_acc_1224_nl[15:0];
  assign nl_Product1_8_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4904:4900]));
  assign Product1_8_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5544:5540]));
  assign Product1_9_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1223_nl = (readslicef_20_16_4(Product1_8_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1223_nl = nl_Accum2_acc_1223_nl[15:0];
  assign nl_Accum2_acc_1232_nl = Accum2_acc_1226_nl + Accum2_acc_1225_nl + Accum2_acc_1224_nl
      + Accum2_acc_1223_nl;
  assign Accum2_acc_1232_nl = nl_Accum2_acc_1232_nl[15:0];
  assign nl_Product1_10_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6184:6180]));
  assign Product1_10_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6824:6820]));
  assign Product1_11_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1222_nl = (readslicef_20_16_4(Product1_10_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1222_nl = nl_Accum2_acc_1222_nl[15:0];
  assign nl_Product1_12_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7464:7460]));
  assign Product1_12_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8104:8100]));
  assign Product1_13_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1221_nl = (readslicef_20_16_4(Product1_12_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1221_nl = nl_Accum2_acc_1221_nl[15:0];
  assign nl_Accum2_acc_1228_nl = Accum2_acc_1222_nl + Accum2_acc_1221_nl;
  assign Accum2_acc_1228_nl = nl_Accum2_acc_1228_nl[15:0];
  assign nl_Accum2_acc_1876_nl = (Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[424:420]);
  assign Accum2_acc_1876_nl = nl_Accum2_acc_1876_nl[9:0];
  assign nl_Product1_1_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[424:420]));
  assign Product1_1_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1227_nl = ({Accum2_acc_1876_nl , (Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1227_nl = nl_Accum2_acc_1227_nl[15:0];
  assign nl_Accum2_acc_1231_nl = Accum2_acc_1228_nl + Accum2_acc_1227_nl;
  assign Accum2_acc_1231_nl = nl_Accum2_acc_1231_nl[15:0];
  assign nl_Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1232_nl + Accum2_acc_1231_nl;
  assign Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1 = (Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1069:1065]));
  assign Product1_2_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1709:1705]));
  assign Product1_3_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1239_nl = (readslicef_20_16_4(Product1_2_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1239_nl = nl_Accum2_acc_1239_nl[15:0];
  assign nl_Product1_4_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2349:2345]));
  assign Product1_4_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2989:2985]));
  assign Product1_5_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1238_nl = (readslicef_20_16_4(Product1_4_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1238_nl = nl_Accum2_acc_1238_nl[15:0];
  assign nl_Product1_6_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3629:3625]));
  assign Product1_6_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4269:4265]));
  assign Product1_7_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1237_nl = (readslicef_20_16_4(Product1_6_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1237_nl = nl_Accum2_acc_1237_nl[15:0];
  assign nl_Product1_8_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4909:4905]));
  assign Product1_8_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5549:5545]));
  assign Product1_9_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1236_nl = (readslicef_20_16_4(Product1_8_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1236_nl = nl_Accum2_acc_1236_nl[15:0];
  assign nl_Accum2_acc_1245_nl = Accum2_acc_1239_nl + Accum2_acc_1238_nl + Accum2_acc_1237_nl
      + Accum2_acc_1236_nl;
  assign Accum2_acc_1245_nl = nl_Accum2_acc_1245_nl[15:0];
  assign nl_Product1_10_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6189:6185]));
  assign Product1_10_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6829:6825]));
  assign Product1_11_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1235_nl = (readslicef_20_16_4(Product1_10_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1235_nl = nl_Accum2_acc_1235_nl[15:0];
  assign nl_Product1_12_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7469:7465]));
  assign Product1_12_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8109:8105]));
  assign Product1_13_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1234_nl = (readslicef_20_16_4(Product1_12_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1234_nl = nl_Accum2_acc_1234_nl[15:0];
  assign nl_Accum2_acc_1241_nl = Accum2_acc_1235_nl + Accum2_acc_1234_nl;
  assign Accum2_acc_1241_nl = nl_Accum2_acc_1241_nl[15:0];
  assign nl_Accum2_acc_1877_nl = (Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[429:425]);
  assign Accum2_acc_1877_nl = nl_Accum2_acc_1877_nl[9:0];
  assign nl_Product1_1_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[429:425]));
  assign Product1_1_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1240_nl = ({Accum2_acc_1877_nl , (Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1240_nl = nl_Accum2_acc_1240_nl[15:0];
  assign nl_Accum2_acc_1244_nl = Accum2_acc_1241_nl + Accum2_acc_1240_nl;
  assign Accum2_acc_1244_nl = nl_Accum2_acc_1244_nl[15:0];
  assign nl_Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1245_nl + Accum2_acc_1244_nl;
  assign Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1 = (Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1074:1070]));
  assign Product1_2_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1714:1710]));
  assign Product1_3_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1252_nl = (readslicef_20_16_4(Product1_2_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1252_nl = nl_Accum2_acc_1252_nl[15:0];
  assign nl_Product1_4_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2354:2350]));
  assign Product1_4_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2994:2990]));
  assign Product1_5_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1251_nl = (readslicef_20_16_4(Product1_4_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1251_nl = nl_Accum2_acc_1251_nl[15:0];
  assign nl_Product1_6_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3634:3630]));
  assign Product1_6_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4274:4270]));
  assign Product1_7_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1250_nl = (readslicef_20_16_4(Product1_6_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1250_nl = nl_Accum2_acc_1250_nl[15:0];
  assign nl_Product1_8_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4914:4910]));
  assign Product1_8_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5554:5550]));
  assign Product1_9_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1249_nl = (readslicef_20_16_4(Product1_8_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1249_nl = nl_Accum2_acc_1249_nl[15:0];
  assign nl_Accum2_acc_1258_nl = Accum2_acc_1252_nl + Accum2_acc_1251_nl + Accum2_acc_1250_nl
      + Accum2_acc_1249_nl;
  assign Accum2_acc_1258_nl = nl_Accum2_acc_1258_nl[15:0];
  assign nl_Product1_10_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6194:6190]));
  assign Product1_10_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6834:6830]));
  assign Product1_11_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1248_nl = (readslicef_20_16_4(Product1_10_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1248_nl = nl_Accum2_acc_1248_nl[15:0];
  assign nl_Product1_12_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7474:7470]));
  assign Product1_12_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8114:8110]));
  assign Product1_13_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1247_nl = (readslicef_20_16_4(Product1_12_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1247_nl = nl_Accum2_acc_1247_nl[15:0];
  assign nl_Accum2_acc_1254_nl = Accum2_acc_1248_nl + Accum2_acc_1247_nl;
  assign Accum2_acc_1254_nl = nl_Accum2_acc_1254_nl[15:0];
  assign nl_Accum2_acc_1878_nl = (Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[434:430]);
  assign Accum2_acc_1878_nl = nl_Accum2_acc_1878_nl[9:0];
  assign nl_Product1_1_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[434:430]));
  assign Product1_1_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1253_nl = ({Accum2_acc_1878_nl , (Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1253_nl = nl_Accum2_acc_1253_nl[15:0];
  assign nl_Accum2_acc_1257_nl = Accum2_acc_1254_nl + Accum2_acc_1253_nl;
  assign Accum2_acc_1257_nl = nl_Accum2_acc_1257_nl[15:0];
  assign nl_Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1258_nl + Accum2_acc_1257_nl;
  assign Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1 = (Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1079:1075]));
  assign Product1_2_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1719:1715]));
  assign Product1_3_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1265_nl = (readslicef_20_16_4(Product1_2_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1265_nl = nl_Accum2_acc_1265_nl[15:0];
  assign nl_Product1_4_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2359:2355]));
  assign Product1_4_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[2999:2995]));
  assign Product1_5_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1264_nl = (readslicef_20_16_4(Product1_4_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1264_nl = nl_Accum2_acc_1264_nl[15:0];
  assign nl_Product1_6_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3639:3635]));
  assign Product1_6_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4279:4275]));
  assign Product1_7_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1263_nl = (readslicef_20_16_4(Product1_6_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1263_nl = nl_Accum2_acc_1263_nl[15:0];
  assign nl_Product1_8_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4919:4915]));
  assign Product1_8_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5559:5555]));
  assign Product1_9_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1262_nl = (readslicef_20_16_4(Product1_8_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1262_nl = nl_Accum2_acc_1262_nl[15:0];
  assign nl_Accum2_acc_1271_nl = Accum2_acc_1265_nl + Accum2_acc_1264_nl + Accum2_acc_1263_nl
      + Accum2_acc_1262_nl;
  assign Accum2_acc_1271_nl = nl_Accum2_acc_1271_nl[15:0];
  assign nl_Product1_10_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6199:6195]));
  assign Product1_10_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6839:6835]));
  assign Product1_11_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1261_nl = (readslicef_20_16_4(Product1_10_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1261_nl = nl_Accum2_acc_1261_nl[15:0];
  assign nl_Product1_12_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7479:7475]));
  assign Product1_12_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8119:8115]));
  assign Product1_13_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1260_nl = (readslicef_20_16_4(Product1_12_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1260_nl = nl_Accum2_acc_1260_nl[15:0];
  assign nl_Accum2_acc_1267_nl = Accum2_acc_1261_nl + Accum2_acc_1260_nl;
  assign Accum2_acc_1267_nl = nl_Accum2_acc_1267_nl[15:0];
  assign nl_Accum2_acc_1879_nl = (Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[439:435]);
  assign Accum2_acc_1879_nl = nl_Accum2_acc_1879_nl[9:0];
  assign nl_Product1_1_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[439:435]));
  assign Product1_1_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1266_nl = ({Accum2_acc_1879_nl , (Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1266_nl = nl_Accum2_acc_1266_nl[15:0];
  assign nl_Accum2_acc_1270_nl = Accum2_acc_1267_nl + Accum2_acc_1266_nl;
  assign Accum2_acc_1270_nl = nl_Accum2_acc_1270_nl[15:0];
  assign nl_Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1271_nl + Accum2_acc_1270_nl;
  assign Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1 = (Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1084:1080]));
  assign Product1_2_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1724:1720]));
  assign Product1_3_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1278_nl = (readslicef_20_16_4(Product1_2_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1278_nl = nl_Accum2_acc_1278_nl[15:0];
  assign nl_Product1_4_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2364:2360]));
  assign Product1_4_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3004:3000]));
  assign Product1_5_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1277_nl = (readslicef_20_16_4(Product1_4_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1277_nl = nl_Accum2_acc_1277_nl[15:0];
  assign nl_Product1_6_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3644:3640]));
  assign Product1_6_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4284:4280]));
  assign Product1_7_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1276_nl = (readslicef_20_16_4(Product1_6_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1276_nl = nl_Accum2_acc_1276_nl[15:0];
  assign nl_Product1_8_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4924:4920]));
  assign Product1_8_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5564:5560]));
  assign Product1_9_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1275_nl = (readslicef_20_16_4(Product1_8_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1275_nl = nl_Accum2_acc_1275_nl[15:0];
  assign nl_Accum2_acc_1284_nl = Accum2_acc_1278_nl + Accum2_acc_1277_nl + Accum2_acc_1276_nl
      + Accum2_acc_1275_nl;
  assign Accum2_acc_1284_nl = nl_Accum2_acc_1284_nl[15:0];
  assign nl_Product1_10_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6204:6200]));
  assign Product1_10_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6844:6840]));
  assign Product1_11_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1274_nl = (readslicef_20_16_4(Product1_10_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1274_nl = nl_Accum2_acc_1274_nl[15:0];
  assign nl_Product1_12_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7484:7480]));
  assign Product1_12_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8124:8120]));
  assign Product1_13_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1273_nl = (readslicef_20_16_4(Product1_12_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1273_nl = nl_Accum2_acc_1273_nl[15:0];
  assign nl_Accum2_acc_1280_nl = Accum2_acc_1274_nl + Accum2_acc_1273_nl;
  assign Accum2_acc_1280_nl = nl_Accum2_acc_1280_nl[15:0];
  assign nl_Accum2_acc_1880_nl = (Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[444:440]);
  assign Accum2_acc_1880_nl = nl_Accum2_acc_1880_nl[9:0];
  assign nl_Product1_1_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[444:440]));
  assign Product1_1_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1279_nl = ({Accum2_acc_1880_nl , (Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1279_nl = nl_Accum2_acc_1279_nl[15:0];
  assign nl_Accum2_acc_1283_nl = Accum2_acc_1280_nl + Accum2_acc_1279_nl;
  assign Accum2_acc_1283_nl = nl_Accum2_acc_1283_nl[15:0];
  assign nl_Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1284_nl + Accum2_acc_1283_nl;
  assign Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1 = (Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1089:1085]));
  assign Product1_2_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1729:1725]));
  assign Product1_3_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1291_nl = (readslicef_20_16_4(Product1_2_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1291_nl = nl_Accum2_acc_1291_nl[15:0];
  assign nl_Product1_4_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2369:2365]));
  assign Product1_4_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3009:3005]));
  assign Product1_5_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1290_nl = (readslicef_20_16_4(Product1_4_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1290_nl = nl_Accum2_acc_1290_nl[15:0];
  assign nl_Product1_6_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3649:3645]));
  assign Product1_6_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4289:4285]));
  assign Product1_7_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1289_nl = (readslicef_20_16_4(Product1_6_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1289_nl = nl_Accum2_acc_1289_nl[15:0];
  assign nl_Product1_8_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4929:4925]));
  assign Product1_8_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5569:5565]));
  assign Product1_9_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1288_nl = (readslicef_20_16_4(Product1_8_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1288_nl = nl_Accum2_acc_1288_nl[15:0];
  assign nl_Accum2_acc_1297_nl = Accum2_acc_1291_nl + Accum2_acc_1290_nl + Accum2_acc_1289_nl
      + Accum2_acc_1288_nl;
  assign Accum2_acc_1297_nl = nl_Accum2_acc_1297_nl[15:0];
  assign nl_Product1_10_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6209:6205]));
  assign Product1_10_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6849:6845]));
  assign Product1_11_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1287_nl = (readslicef_20_16_4(Product1_10_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1287_nl = nl_Accum2_acc_1287_nl[15:0];
  assign nl_Product1_12_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7489:7485]));
  assign Product1_12_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8129:8125]));
  assign Product1_13_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1286_nl = (readslicef_20_16_4(Product1_12_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1286_nl = nl_Accum2_acc_1286_nl[15:0];
  assign nl_Accum2_acc_1293_nl = Accum2_acc_1287_nl + Accum2_acc_1286_nl;
  assign Accum2_acc_1293_nl = nl_Accum2_acc_1293_nl[15:0];
  assign nl_Accum2_acc_1881_nl = (Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[449:445]);
  assign Accum2_acc_1881_nl = nl_Accum2_acc_1881_nl[9:0];
  assign nl_Product1_1_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[449:445]));
  assign Product1_1_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1292_nl = ({Accum2_acc_1881_nl , (Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1292_nl = nl_Accum2_acc_1292_nl[15:0];
  assign nl_Accum2_acc_1296_nl = Accum2_acc_1293_nl + Accum2_acc_1292_nl;
  assign Accum2_acc_1296_nl = nl_Accum2_acc_1296_nl[15:0];
  assign nl_Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1297_nl + Accum2_acc_1296_nl;
  assign Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1 = (Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1094:1090]));
  assign Product1_2_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1734:1730]));
  assign Product1_3_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1304_nl = (readslicef_20_16_4(Product1_2_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1304_nl = nl_Accum2_acc_1304_nl[15:0];
  assign nl_Product1_4_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2374:2370]));
  assign Product1_4_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3014:3010]));
  assign Product1_5_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1303_nl = (readslicef_20_16_4(Product1_4_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1303_nl = nl_Accum2_acc_1303_nl[15:0];
  assign nl_Product1_6_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3654:3650]));
  assign Product1_6_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4294:4290]));
  assign Product1_7_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1302_nl = (readslicef_20_16_4(Product1_6_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1302_nl = nl_Accum2_acc_1302_nl[15:0];
  assign nl_Product1_8_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4934:4930]));
  assign Product1_8_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5574:5570]));
  assign Product1_9_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1301_nl = (readslicef_20_16_4(Product1_8_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1301_nl = nl_Accum2_acc_1301_nl[15:0];
  assign nl_Accum2_acc_1310_nl = Accum2_acc_1304_nl + Accum2_acc_1303_nl + Accum2_acc_1302_nl
      + Accum2_acc_1301_nl;
  assign Accum2_acc_1310_nl = nl_Accum2_acc_1310_nl[15:0];
  assign nl_Product1_10_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6214:6210]));
  assign Product1_10_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6854:6850]));
  assign Product1_11_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1300_nl = (readslicef_20_16_4(Product1_10_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1300_nl = nl_Accum2_acc_1300_nl[15:0];
  assign nl_Product1_12_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7494:7490]));
  assign Product1_12_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8134:8130]));
  assign Product1_13_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1299_nl = (readslicef_20_16_4(Product1_12_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1299_nl = nl_Accum2_acc_1299_nl[15:0];
  assign nl_Accum2_acc_1306_nl = Accum2_acc_1300_nl + Accum2_acc_1299_nl;
  assign Accum2_acc_1306_nl = nl_Accum2_acc_1306_nl[15:0];
  assign nl_Accum2_acc_1882_nl = (Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[454:450]);
  assign Accum2_acc_1882_nl = nl_Accum2_acc_1882_nl[9:0];
  assign nl_Product1_1_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[454:450]));
  assign Product1_1_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1305_nl = ({Accum2_acc_1882_nl , (Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1305_nl = nl_Accum2_acc_1305_nl[15:0];
  assign nl_Accum2_acc_1309_nl = Accum2_acc_1306_nl + Accum2_acc_1305_nl;
  assign Accum2_acc_1309_nl = nl_Accum2_acc_1309_nl[15:0];
  assign nl_Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1310_nl + Accum2_acc_1309_nl;
  assign Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1 = (Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1099:1095]));
  assign Product1_2_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1739:1735]));
  assign Product1_3_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1317_nl = (readslicef_20_16_4(Product1_2_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1317_nl = nl_Accum2_acc_1317_nl[15:0];
  assign nl_Product1_4_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2379:2375]));
  assign Product1_4_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3019:3015]));
  assign Product1_5_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1316_nl = (readslicef_20_16_4(Product1_4_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1316_nl = nl_Accum2_acc_1316_nl[15:0];
  assign nl_Product1_6_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3659:3655]));
  assign Product1_6_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4299:4295]));
  assign Product1_7_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1315_nl = (readslicef_20_16_4(Product1_6_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1315_nl = nl_Accum2_acc_1315_nl[15:0];
  assign nl_Product1_8_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4939:4935]));
  assign Product1_8_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5579:5575]));
  assign Product1_9_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1314_nl = (readslicef_20_16_4(Product1_8_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1314_nl = nl_Accum2_acc_1314_nl[15:0];
  assign nl_Accum2_acc_1323_nl = Accum2_acc_1317_nl + Accum2_acc_1316_nl + Accum2_acc_1315_nl
      + Accum2_acc_1314_nl;
  assign Accum2_acc_1323_nl = nl_Accum2_acc_1323_nl[15:0];
  assign nl_Product1_10_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6219:6215]));
  assign Product1_10_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6859:6855]));
  assign Product1_11_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1313_nl = (readslicef_20_16_4(Product1_10_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1313_nl = nl_Accum2_acc_1313_nl[15:0];
  assign nl_Product1_12_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7499:7495]));
  assign Product1_12_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8139:8135]));
  assign Product1_13_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1312_nl = (readslicef_20_16_4(Product1_12_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1312_nl = nl_Accum2_acc_1312_nl[15:0];
  assign nl_Accum2_acc_1319_nl = Accum2_acc_1313_nl + Accum2_acc_1312_nl;
  assign Accum2_acc_1319_nl = nl_Accum2_acc_1319_nl[15:0];
  assign nl_Accum2_acc_1883_nl = (Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[459:455]);
  assign Accum2_acc_1883_nl = nl_Accum2_acc_1883_nl[9:0];
  assign nl_Product1_1_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[459:455]));
  assign Product1_1_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1318_nl = ({Accum2_acc_1883_nl , (Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1318_nl = nl_Accum2_acc_1318_nl[15:0];
  assign nl_Accum2_acc_1322_nl = Accum2_acc_1319_nl + Accum2_acc_1318_nl;
  assign Accum2_acc_1322_nl = nl_Accum2_acc_1322_nl[15:0];
  assign nl_Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1323_nl + Accum2_acc_1322_nl;
  assign Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1 = (Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1104:1100]));
  assign Product1_2_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1744:1740]));
  assign Product1_3_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1330_nl = (readslicef_20_16_4(Product1_2_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1330_nl = nl_Accum2_acc_1330_nl[15:0];
  assign nl_Product1_4_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2384:2380]));
  assign Product1_4_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3024:3020]));
  assign Product1_5_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1329_nl = (readslicef_20_16_4(Product1_4_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1329_nl = nl_Accum2_acc_1329_nl[15:0];
  assign nl_Product1_6_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3664:3660]));
  assign Product1_6_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4304:4300]));
  assign Product1_7_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1328_nl = (readslicef_20_16_4(Product1_6_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1328_nl = nl_Accum2_acc_1328_nl[15:0];
  assign nl_Product1_8_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4944:4940]));
  assign Product1_8_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5584:5580]));
  assign Product1_9_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1327_nl = (readslicef_20_16_4(Product1_8_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1327_nl = nl_Accum2_acc_1327_nl[15:0];
  assign nl_Accum2_acc_1336_nl = Accum2_acc_1330_nl + Accum2_acc_1329_nl + Accum2_acc_1328_nl
      + Accum2_acc_1327_nl;
  assign Accum2_acc_1336_nl = nl_Accum2_acc_1336_nl[15:0];
  assign nl_Product1_10_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6224:6220]));
  assign Product1_10_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6864:6860]));
  assign Product1_11_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1326_nl = (readslicef_20_16_4(Product1_10_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1326_nl = nl_Accum2_acc_1326_nl[15:0];
  assign nl_Product1_12_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7504:7500]));
  assign Product1_12_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8144:8140]));
  assign Product1_13_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1325_nl = (readslicef_20_16_4(Product1_12_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1325_nl = nl_Accum2_acc_1325_nl[15:0];
  assign nl_Accum2_acc_1332_nl = Accum2_acc_1326_nl + Accum2_acc_1325_nl;
  assign Accum2_acc_1332_nl = nl_Accum2_acc_1332_nl[15:0];
  assign nl_Accum2_acc_1884_nl = (Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[464:460]);
  assign Accum2_acc_1884_nl = nl_Accum2_acc_1884_nl[9:0];
  assign nl_Product1_1_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[464:460]));
  assign Product1_1_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1331_nl = ({Accum2_acc_1884_nl , (Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1331_nl = nl_Accum2_acc_1331_nl[15:0];
  assign nl_Accum2_acc_1335_nl = Accum2_acc_1332_nl + Accum2_acc_1331_nl;
  assign Accum2_acc_1335_nl = nl_Accum2_acc_1335_nl[15:0];
  assign nl_Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1336_nl + Accum2_acc_1335_nl;
  assign Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1 = (Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1109:1105]));
  assign Product1_2_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1749:1745]));
  assign Product1_3_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1343_nl = (readslicef_20_16_4(Product1_2_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1343_nl = nl_Accum2_acc_1343_nl[15:0];
  assign nl_Product1_4_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2389:2385]));
  assign Product1_4_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3029:3025]));
  assign Product1_5_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1342_nl = (readslicef_20_16_4(Product1_4_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1342_nl = nl_Accum2_acc_1342_nl[15:0];
  assign nl_Product1_6_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3669:3665]));
  assign Product1_6_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4309:4305]));
  assign Product1_7_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1341_nl = (readslicef_20_16_4(Product1_6_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1341_nl = nl_Accum2_acc_1341_nl[15:0];
  assign nl_Product1_8_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4949:4945]));
  assign Product1_8_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5589:5585]));
  assign Product1_9_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1340_nl = (readslicef_20_16_4(Product1_8_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1340_nl = nl_Accum2_acc_1340_nl[15:0];
  assign nl_Accum2_acc_1349_nl = Accum2_acc_1343_nl + Accum2_acc_1342_nl + Accum2_acc_1341_nl
      + Accum2_acc_1340_nl;
  assign Accum2_acc_1349_nl = nl_Accum2_acc_1349_nl[15:0];
  assign nl_Product1_10_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6229:6225]));
  assign Product1_10_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6869:6865]));
  assign Product1_11_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1339_nl = (readslicef_20_16_4(Product1_10_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1339_nl = nl_Accum2_acc_1339_nl[15:0];
  assign nl_Product1_12_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7509:7505]));
  assign Product1_12_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8149:8145]));
  assign Product1_13_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1338_nl = (readslicef_20_16_4(Product1_12_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1338_nl = nl_Accum2_acc_1338_nl[15:0];
  assign nl_Accum2_acc_1345_nl = Accum2_acc_1339_nl + Accum2_acc_1338_nl;
  assign Accum2_acc_1345_nl = nl_Accum2_acc_1345_nl[15:0];
  assign nl_Accum2_acc_1885_nl = (Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[469:465]);
  assign Accum2_acc_1885_nl = nl_Accum2_acc_1885_nl[9:0];
  assign nl_Product1_1_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[469:465]));
  assign Product1_1_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1344_nl = ({Accum2_acc_1885_nl , (Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1344_nl = nl_Accum2_acc_1344_nl[15:0];
  assign nl_Accum2_acc_1348_nl = Accum2_acc_1345_nl + Accum2_acc_1344_nl;
  assign Accum2_acc_1348_nl = nl_Accum2_acc_1348_nl[15:0];
  assign nl_Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1349_nl + Accum2_acc_1348_nl;
  assign Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1 = (Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1114:1110]));
  assign Product1_2_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1754:1750]));
  assign Product1_3_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1356_nl = (readslicef_20_16_4(Product1_2_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1356_nl = nl_Accum2_acc_1356_nl[15:0];
  assign nl_Product1_4_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2394:2390]));
  assign Product1_4_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3034:3030]));
  assign Product1_5_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1355_nl = (readslicef_20_16_4(Product1_4_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1355_nl = nl_Accum2_acc_1355_nl[15:0];
  assign nl_Product1_6_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3674:3670]));
  assign Product1_6_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4314:4310]));
  assign Product1_7_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1354_nl = (readslicef_20_16_4(Product1_6_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1354_nl = nl_Accum2_acc_1354_nl[15:0];
  assign nl_Product1_8_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4954:4950]));
  assign Product1_8_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5594:5590]));
  assign Product1_9_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1353_nl = (readslicef_20_16_4(Product1_8_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1353_nl = nl_Accum2_acc_1353_nl[15:0];
  assign nl_Accum2_acc_1362_nl = Accum2_acc_1356_nl + Accum2_acc_1355_nl + Accum2_acc_1354_nl
      + Accum2_acc_1353_nl;
  assign Accum2_acc_1362_nl = nl_Accum2_acc_1362_nl[15:0];
  assign nl_Product1_10_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6234:6230]));
  assign Product1_10_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6874:6870]));
  assign Product1_11_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1352_nl = (readslicef_20_16_4(Product1_10_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1352_nl = nl_Accum2_acc_1352_nl[15:0];
  assign nl_Product1_12_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7514:7510]));
  assign Product1_12_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8154:8150]));
  assign Product1_13_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1351_nl = (readslicef_20_16_4(Product1_12_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1351_nl = nl_Accum2_acc_1351_nl[15:0];
  assign nl_Accum2_acc_1358_nl = Accum2_acc_1352_nl + Accum2_acc_1351_nl;
  assign Accum2_acc_1358_nl = nl_Accum2_acc_1358_nl[15:0];
  assign nl_Accum2_acc_1886_nl = (Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[474:470]);
  assign Accum2_acc_1886_nl = nl_Accum2_acc_1886_nl[9:0];
  assign nl_Product1_1_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[474:470]));
  assign Product1_1_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1357_nl = ({Accum2_acc_1886_nl , (Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1357_nl = nl_Accum2_acc_1357_nl[15:0];
  assign nl_Accum2_acc_1361_nl = Accum2_acc_1358_nl + Accum2_acc_1357_nl;
  assign Accum2_acc_1361_nl = nl_Accum2_acc_1361_nl[15:0];
  assign nl_Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1362_nl + Accum2_acc_1361_nl;
  assign Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1 = (Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1119:1115]));
  assign Product1_2_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1759:1755]));
  assign Product1_3_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1369_nl = (readslicef_20_16_4(Product1_2_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1369_nl = nl_Accum2_acc_1369_nl[15:0];
  assign nl_Product1_4_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2399:2395]));
  assign Product1_4_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3039:3035]));
  assign Product1_5_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1368_nl = (readslicef_20_16_4(Product1_4_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1368_nl = nl_Accum2_acc_1368_nl[15:0];
  assign nl_Product1_6_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3679:3675]));
  assign Product1_6_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4319:4315]));
  assign Product1_7_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1367_nl = (readslicef_20_16_4(Product1_6_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1367_nl = nl_Accum2_acc_1367_nl[15:0];
  assign nl_Product1_8_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4959:4955]));
  assign Product1_8_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5599:5595]));
  assign Product1_9_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1366_nl = (readslicef_20_16_4(Product1_8_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1366_nl = nl_Accum2_acc_1366_nl[15:0];
  assign nl_Accum2_acc_1375_nl = Accum2_acc_1369_nl + Accum2_acc_1368_nl + Accum2_acc_1367_nl
      + Accum2_acc_1366_nl;
  assign Accum2_acc_1375_nl = nl_Accum2_acc_1375_nl[15:0];
  assign nl_Product1_10_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6239:6235]));
  assign Product1_10_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6879:6875]));
  assign Product1_11_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1365_nl = (readslicef_20_16_4(Product1_10_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1365_nl = nl_Accum2_acc_1365_nl[15:0];
  assign nl_Product1_12_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7519:7515]));
  assign Product1_12_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8159:8155]));
  assign Product1_13_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1364_nl = (readslicef_20_16_4(Product1_12_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1364_nl = nl_Accum2_acc_1364_nl[15:0];
  assign nl_Accum2_acc_1371_nl = Accum2_acc_1365_nl + Accum2_acc_1364_nl;
  assign Accum2_acc_1371_nl = nl_Accum2_acc_1371_nl[15:0];
  assign nl_Accum2_acc_1887_nl = (Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[479:475]);
  assign Accum2_acc_1887_nl = nl_Accum2_acc_1887_nl[9:0];
  assign nl_Product1_1_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[479:475]));
  assign Product1_1_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1370_nl = ({Accum2_acc_1887_nl , (Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1370_nl = nl_Accum2_acc_1370_nl[15:0];
  assign nl_Accum2_acc_1374_nl = Accum2_acc_1371_nl + Accum2_acc_1370_nl;
  assign Accum2_acc_1374_nl = nl_Accum2_acc_1374_nl[15:0];
  assign nl_Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1375_nl + Accum2_acc_1374_nl;
  assign Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1 = (Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1124:1120]));
  assign Product1_2_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1764:1760]));
  assign Product1_3_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1382_nl = (readslicef_20_16_4(Product1_2_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1382_nl = nl_Accum2_acc_1382_nl[15:0];
  assign nl_Product1_4_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2404:2400]));
  assign Product1_4_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3044:3040]));
  assign Product1_5_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1381_nl = (readslicef_20_16_4(Product1_4_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1381_nl = nl_Accum2_acc_1381_nl[15:0];
  assign nl_Product1_6_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3684:3680]));
  assign Product1_6_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4324:4320]));
  assign Product1_7_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1380_nl = (readslicef_20_16_4(Product1_6_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1380_nl = nl_Accum2_acc_1380_nl[15:0];
  assign nl_Product1_8_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4964:4960]));
  assign Product1_8_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5604:5600]));
  assign Product1_9_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1379_nl = (readslicef_20_16_4(Product1_8_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1379_nl = nl_Accum2_acc_1379_nl[15:0];
  assign nl_Accum2_acc_1388_nl = Accum2_acc_1382_nl + Accum2_acc_1381_nl + Accum2_acc_1380_nl
      + Accum2_acc_1379_nl;
  assign Accum2_acc_1388_nl = nl_Accum2_acc_1388_nl[15:0];
  assign nl_Product1_10_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6244:6240]));
  assign Product1_10_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6884:6880]));
  assign Product1_11_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1378_nl = (readslicef_20_16_4(Product1_10_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1378_nl = nl_Accum2_acc_1378_nl[15:0];
  assign nl_Product1_12_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7524:7520]));
  assign Product1_12_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8164:8160]));
  assign Product1_13_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1377_nl = (readslicef_20_16_4(Product1_12_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1377_nl = nl_Accum2_acc_1377_nl[15:0];
  assign nl_Accum2_acc_1384_nl = Accum2_acc_1378_nl + Accum2_acc_1377_nl;
  assign Accum2_acc_1384_nl = nl_Accum2_acc_1384_nl[15:0];
  assign nl_Accum2_acc_1888_nl = (Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[484:480]);
  assign Accum2_acc_1888_nl = nl_Accum2_acc_1888_nl[9:0];
  assign nl_Product1_1_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[484:480]));
  assign Product1_1_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1383_nl = ({Accum2_acc_1888_nl , (Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1383_nl = nl_Accum2_acc_1383_nl[15:0];
  assign nl_Accum2_acc_1387_nl = Accum2_acc_1384_nl + Accum2_acc_1383_nl;
  assign Accum2_acc_1387_nl = nl_Accum2_acc_1387_nl[15:0];
  assign nl_Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1388_nl + Accum2_acc_1387_nl;
  assign Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1 = (Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1129:1125]));
  assign Product1_2_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1769:1765]));
  assign Product1_3_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1395_nl = (readslicef_20_16_4(Product1_2_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1395_nl = nl_Accum2_acc_1395_nl[15:0];
  assign nl_Product1_4_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2409:2405]));
  assign Product1_4_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3049:3045]));
  assign Product1_5_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1394_nl = (readslicef_20_16_4(Product1_4_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1394_nl = nl_Accum2_acc_1394_nl[15:0];
  assign nl_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3689:3685]));
  assign Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4329:4325]));
  assign Product1_7_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1393_nl = (readslicef_20_16_4(Product1_6_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1393_nl = nl_Accum2_acc_1393_nl[15:0];
  assign nl_Product1_8_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4969:4965]));
  assign Product1_8_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5609:5605]));
  assign Product1_9_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1392_nl = (readslicef_20_16_4(Product1_8_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1392_nl = nl_Accum2_acc_1392_nl[15:0];
  assign nl_Accum2_acc_1401_nl = Accum2_acc_1395_nl + Accum2_acc_1394_nl + Accum2_acc_1393_nl
      + Accum2_acc_1392_nl;
  assign Accum2_acc_1401_nl = nl_Accum2_acc_1401_nl[15:0];
  assign nl_Product1_10_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6249:6245]));
  assign Product1_10_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6889:6885]));
  assign Product1_11_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1391_nl = (readslicef_20_16_4(Product1_10_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1391_nl = nl_Accum2_acc_1391_nl[15:0];
  assign nl_Product1_12_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7529:7525]));
  assign Product1_12_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8169:8165]));
  assign Product1_13_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1390_nl = (readslicef_20_16_4(Product1_12_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1390_nl = nl_Accum2_acc_1390_nl[15:0];
  assign nl_Accum2_acc_1397_nl = Accum2_acc_1391_nl + Accum2_acc_1390_nl;
  assign Accum2_acc_1397_nl = nl_Accum2_acc_1397_nl[15:0];
  assign nl_Accum2_acc_1889_nl = (Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[489:485]);
  assign Accum2_acc_1889_nl = nl_Accum2_acc_1889_nl[9:0];
  assign nl_Product1_1_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[489:485]));
  assign Product1_1_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1396_nl = ({Accum2_acc_1889_nl , (Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1396_nl = nl_Accum2_acc_1396_nl[15:0];
  assign nl_Accum2_acc_1400_nl = Accum2_acc_1397_nl + Accum2_acc_1396_nl;
  assign Accum2_acc_1400_nl = nl_Accum2_acc_1400_nl[15:0];
  assign nl_Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1401_nl + Accum2_acc_1400_nl;
  assign Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1 = (Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1134:1130]));
  assign Product1_2_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1774:1770]));
  assign Product1_3_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1408_nl = (readslicef_20_16_4(Product1_2_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1408_nl = nl_Accum2_acc_1408_nl[15:0];
  assign nl_Product1_4_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2414:2410]));
  assign Product1_4_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3054:3050]));
  assign Product1_5_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1407_nl = (readslicef_20_16_4(Product1_4_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1407_nl = nl_Accum2_acc_1407_nl[15:0];
  assign nl_Product1_6_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3694:3690]));
  assign Product1_6_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4334:4330]));
  assign Product1_7_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1406_nl = (readslicef_20_16_4(Product1_6_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1406_nl = nl_Accum2_acc_1406_nl[15:0];
  assign nl_Product1_8_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4974:4970]));
  assign Product1_8_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5614:5610]));
  assign Product1_9_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1405_nl = (readslicef_20_16_4(Product1_8_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1405_nl = nl_Accum2_acc_1405_nl[15:0];
  assign nl_Accum2_acc_1414_nl = Accum2_acc_1408_nl + Accum2_acc_1407_nl + Accum2_acc_1406_nl
      + Accum2_acc_1405_nl;
  assign Accum2_acc_1414_nl = nl_Accum2_acc_1414_nl[15:0];
  assign nl_Product1_10_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6254:6250]));
  assign Product1_10_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6894:6890]));
  assign Product1_11_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1404_nl = (readslicef_20_16_4(Product1_10_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1404_nl = nl_Accum2_acc_1404_nl[15:0];
  assign nl_Product1_12_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7534:7530]));
  assign Product1_12_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8174:8170]));
  assign Product1_13_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1403_nl = (readslicef_20_16_4(Product1_12_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1403_nl = nl_Accum2_acc_1403_nl[15:0];
  assign nl_Accum2_acc_1410_nl = Accum2_acc_1404_nl + Accum2_acc_1403_nl;
  assign Accum2_acc_1410_nl = nl_Accum2_acc_1410_nl[15:0];
  assign nl_Accum2_acc_1890_nl = (Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[494:490]);
  assign Accum2_acc_1890_nl = nl_Accum2_acc_1890_nl[9:0];
  assign nl_Product1_1_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[494:490]));
  assign Product1_1_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1409_nl = ({Accum2_acc_1890_nl , (Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1409_nl = nl_Accum2_acc_1409_nl[15:0];
  assign nl_Accum2_acc_1413_nl = Accum2_acc_1410_nl + Accum2_acc_1409_nl;
  assign Accum2_acc_1413_nl = nl_Accum2_acc_1413_nl[15:0];
  assign nl_Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1414_nl + Accum2_acc_1413_nl;
  assign Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1 = (Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1139:1135]));
  assign Product1_2_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1779:1775]));
  assign Product1_3_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1421_nl = (readslicef_20_16_4(Product1_2_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1421_nl = nl_Accum2_acc_1421_nl[15:0];
  assign nl_Product1_4_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2419:2415]));
  assign Product1_4_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3059:3055]));
  assign Product1_5_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1420_nl = (readslicef_20_16_4(Product1_4_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1420_nl = nl_Accum2_acc_1420_nl[15:0];
  assign nl_Product1_6_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3699:3695]));
  assign Product1_6_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4339:4335]));
  assign Product1_7_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1419_nl = (readslicef_20_16_4(Product1_6_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1419_nl = nl_Accum2_acc_1419_nl[15:0];
  assign nl_Product1_8_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4979:4975]));
  assign Product1_8_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5619:5615]));
  assign Product1_9_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1418_nl = (readslicef_20_16_4(Product1_8_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1418_nl = nl_Accum2_acc_1418_nl[15:0];
  assign nl_Accum2_acc_1427_nl = Accum2_acc_1421_nl + Accum2_acc_1420_nl + Accum2_acc_1419_nl
      + Accum2_acc_1418_nl;
  assign Accum2_acc_1427_nl = nl_Accum2_acc_1427_nl[15:0];
  assign nl_Product1_10_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6259:6255]));
  assign Product1_10_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6899:6895]));
  assign Product1_11_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1417_nl = (readslicef_20_16_4(Product1_10_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1417_nl = nl_Accum2_acc_1417_nl[15:0];
  assign nl_Product1_12_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7539:7535]));
  assign Product1_12_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8179:8175]));
  assign Product1_13_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1416_nl = (readslicef_20_16_4(Product1_12_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1416_nl = nl_Accum2_acc_1416_nl[15:0];
  assign nl_Accum2_acc_1423_nl = Accum2_acc_1417_nl + Accum2_acc_1416_nl;
  assign Accum2_acc_1423_nl = nl_Accum2_acc_1423_nl[15:0];
  assign nl_Accum2_acc_1891_nl = (Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[499:495]);
  assign Accum2_acc_1891_nl = nl_Accum2_acc_1891_nl[9:0];
  assign nl_Product1_1_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[499:495]));
  assign Product1_1_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1422_nl = ({Accum2_acc_1891_nl , (Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1422_nl = nl_Accum2_acc_1422_nl[15:0];
  assign nl_Accum2_acc_1426_nl = Accum2_acc_1423_nl + Accum2_acc_1422_nl;
  assign Accum2_acc_1426_nl = nl_Accum2_acc_1426_nl[15:0];
  assign nl_Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1427_nl + Accum2_acc_1426_nl;
  assign Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1 = (Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1144:1140]));
  assign Product1_2_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1784:1780]));
  assign Product1_3_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1434_nl = (readslicef_20_16_4(Product1_2_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1434_nl = nl_Accum2_acc_1434_nl[15:0];
  assign nl_Product1_4_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2424:2420]));
  assign Product1_4_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3064:3060]));
  assign Product1_5_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1433_nl = (readslicef_20_16_4(Product1_4_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1433_nl = nl_Accum2_acc_1433_nl[15:0];
  assign nl_Product1_6_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3704:3700]));
  assign Product1_6_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4344:4340]));
  assign Product1_7_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1432_nl = (readslicef_20_16_4(Product1_6_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1432_nl = nl_Accum2_acc_1432_nl[15:0];
  assign nl_Product1_8_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4984:4980]));
  assign Product1_8_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5624:5620]));
  assign Product1_9_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1431_nl = (readslicef_20_16_4(Product1_8_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1431_nl = nl_Accum2_acc_1431_nl[15:0];
  assign nl_Accum2_acc_1440_nl = Accum2_acc_1434_nl + Accum2_acc_1433_nl + Accum2_acc_1432_nl
      + Accum2_acc_1431_nl;
  assign Accum2_acc_1440_nl = nl_Accum2_acc_1440_nl[15:0];
  assign nl_Product1_10_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6264:6260]));
  assign Product1_10_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6904:6900]));
  assign Product1_11_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1430_nl = (readslicef_20_16_4(Product1_10_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1430_nl = nl_Accum2_acc_1430_nl[15:0];
  assign nl_Product1_12_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7544:7540]));
  assign Product1_12_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8184:8180]));
  assign Product1_13_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1429_nl = (readslicef_20_16_4(Product1_12_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1429_nl = nl_Accum2_acc_1429_nl[15:0];
  assign nl_Accum2_acc_1436_nl = Accum2_acc_1430_nl + Accum2_acc_1429_nl;
  assign Accum2_acc_1436_nl = nl_Accum2_acc_1436_nl[15:0];
  assign nl_Accum2_acc_1892_nl = (Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[504:500]);
  assign Accum2_acc_1892_nl = nl_Accum2_acc_1892_nl[9:0];
  assign nl_Product1_1_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[504:500]));
  assign Product1_1_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1435_nl = ({Accum2_acc_1892_nl , (Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1435_nl = nl_Accum2_acc_1435_nl[15:0];
  assign nl_Accum2_acc_1439_nl = Accum2_acc_1436_nl + Accum2_acc_1435_nl;
  assign Accum2_acc_1439_nl = nl_Accum2_acc_1439_nl[15:0];
  assign nl_Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1440_nl + Accum2_acc_1439_nl;
  assign Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1 = (Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1149:1145]));
  assign Product1_2_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1789:1785]));
  assign Product1_3_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1447_nl = (readslicef_20_16_4(Product1_2_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1447_nl = nl_Accum2_acc_1447_nl[15:0];
  assign nl_Product1_4_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2429:2425]));
  assign Product1_4_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3069:3065]));
  assign Product1_5_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1446_nl = (readslicef_20_16_4(Product1_4_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1446_nl = nl_Accum2_acc_1446_nl[15:0];
  assign nl_Product1_6_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3709:3705]));
  assign Product1_6_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4349:4345]));
  assign Product1_7_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1445_nl = (readslicef_20_16_4(Product1_6_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1445_nl = nl_Accum2_acc_1445_nl[15:0];
  assign nl_Product1_8_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4989:4985]));
  assign Product1_8_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5629:5625]));
  assign Product1_9_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1444_nl = (readslicef_20_16_4(Product1_8_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1444_nl = nl_Accum2_acc_1444_nl[15:0];
  assign nl_Accum2_acc_1453_nl = Accum2_acc_1447_nl + Accum2_acc_1446_nl + Accum2_acc_1445_nl
      + Accum2_acc_1444_nl;
  assign Accum2_acc_1453_nl = nl_Accum2_acc_1453_nl[15:0];
  assign nl_Product1_10_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6269:6265]));
  assign Product1_10_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6909:6905]));
  assign Product1_11_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1443_nl = (readslicef_20_16_4(Product1_10_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1443_nl = nl_Accum2_acc_1443_nl[15:0];
  assign nl_Product1_12_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7549:7545]));
  assign Product1_12_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8189:8185]));
  assign Product1_13_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1442_nl = (readslicef_20_16_4(Product1_12_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1442_nl = nl_Accum2_acc_1442_nl[15:0];
  assign nl_Accum2_acc_1449_nl = Accum2_acc_1443_nl + Accum2_acc_1442_nl;
  assign Accum2_acc_1449_nl = nl_Accum2_acc_1449_nl[15:0];
  assign nl_Accum2_acc_1893_nl = (Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[509:505]);
  assign Accum2_acc_1893_nl = nl_Accum2_acc_1893_nl[9:0];
  assign nl_Product1_1_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[509:505]));
  assign Product1_1_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1448_nl = ({Accum2_acc_1893_nl , (Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1448_nl = nl_Accum2_acc_1448_nl[15:0];
  assign nl_Accum2_acc_1452_nl = Accum2_acc_1449_nl + Accum2_acc_1448_nl;
  assign Accum2_acc_1452_nl = nl_Accum2_acc_1452_nl[15:0];
  assign nl_Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1453_nl + Accum2_acc_1452_nl;
  assign Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1 = (Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1154:1150]));
  assign Product1_2_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1794:1790]));
  assign Product1_3_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1460_nl = (readslicef_20_16_4(Product1_2_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1460_nl = nl_Accum2_acc_1460_nl[15:0];
  assign nl_Product1_4_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2434:2430]));
  assign Product1_4_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3074:3070]));
  assign Product1_5_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1459_nl = (readslicef_20_16_4(Product1_4_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1459_nl = nl_Accum2_acc_1459_nl[15:0];
  assign nl_Product1_6_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3714:3710]));
  assign Product1_6_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4354:4350]));
  assign Product1_7_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1458_nl = (readslicef_20_16_4(Product1_6_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1458_nl = nl_Accum2_acc_1458_nl[15:0];
  assign nl_Product1_8_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4994:4990]));
  assign Product1_8_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5634:5630]));
  assign Product1_9_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1457_nl = (readslicef_20_16_4(Product1_8_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1457_nl = nl_Accum2_acc_1457_nl[15:0];
  assign nl_Accum2_acc_1466_nl = Accum2_acc_1460_nl + Accum2_acc_1459_nl + Accum2_acc_1458_nl
      + Accum2_acc_1457_nl;
  assign Accum2_acc_1466_nl = nl_Accum2_acc_1466_nl[15:0];
  assign nl_Product1_10_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6274:6270]));
  assign Product1_10_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6914:6910]));
  assign Product1_11_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1456_nl = (readslicef_20_16_4(Product1_10_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1456_nl = nl_Accum2_acc_1456_nl[15:0];
  assign nl_Product1_12_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7554:7550]));
  assign Product1_12_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8194:8190]));
  assign Product1_13_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1455_nl = (readslicef_20_16_4(Product1_12_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1455_nl = nl_Accum2_acc_1455_nl[15:0];
  assign nl_Accum2_acc_1462_nl = Accum2_acc_1456_nl + Accum2_acc_1455_nl;
  assign Accum2_acc_1462_nl = nl_Accum2_acc_1462_nl[15:0];
  assign nl_Accum2_acc_1894_nl = (Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[514:510]);
  assign Accum2_acc_1894_nl = nl_Accum2_acc_1894_nl[9:0];
  assign nl_Product1_1_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[514:510]));
  assign Product1_1_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1461_nl = ({Accum2_acc_1894_nl , (Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1461_nl = nl_Accum2_acc_1461_nl[15:0];
  assign nl_Accum2_acc_1465_nl = Accum2_acc_1462_nl + Accum2_acc_1461_nl;
  assign Accum2_acc_1465_nl = nl_Accum2_acc_1465_nl[15:0];
  assign nl_Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1466_nl + Accum2_acc_1465_nl;
  assign Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1 = (Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1159:1155]));
  assign Product1_2_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1799:1795]));
  assign Product1_3_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1473_nl = (readslicef_20_16_4(Product1_2_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1473_nl = nl_Accum2_acc_1473_nl[15:0];
  assign nl_Product1_4_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2439:2435]));
  assign Product1_4_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3079:3075]));
  assign Product1_5_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1472_nl = (readslicef_20_16_4(Product1_4_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1472_nl = nl_Accum2_acc_1472_nl[15:0];
  assign nl_Product1_6_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3719:3715]));
  assign Product1_6_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4359:4355]));
  assign Product1_7_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1471_nl = (readslicef_20_16_4(Product1_6_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1471_nl = nl_Accum2_acc_1471_nl[15:0];
  assign nl_Product1_8_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[4999:4995]));
  assign Product1_8_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5639:5635]));
  assign Product1_9_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1470_nl = (readslicef_20_16_4(Product1_8_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1470_nl = nl_Accum2_acc_1470_nl[15:0];
  assign nl_Accum2_acc_1479_nl = Accum2_acc_1473_nl + Accum2_acc_1472_nl + Accum2_acc_1471_nl
      + Accum2_acc_1470_nl;
  assign Accum2_acc_1479_nl = nl_Accum2_acc_1479_nl[15:0];
  assign nl_Product1_10_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6279:6275]));
  assign Product1_10_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6919:6915]));
  assign Product1_11_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1469_nl = (readslicef_20_16_4(Product1_10_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1469_nl = nl_Accum2_acc_1469_nl[15:0];
  assign nl_Product1_12_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7559:7555]));
  assign Product1_12_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8199:8195]));
  assign Product1_13_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1468_nl = (readslicef_20_16_4(Product1_12_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1468_nl = nl_Accum2_acc_1468_nl[15:0];
  assign nl_Accum2_acc_1475_nl = Accum2_acc_1469_nl + Accum2_acc_1468_nl;
  assign Accum2_acc_1475_nl = nl_Accum2_acc_1475_nl[15:0];
  assign nl_Accum2_acc_1895_nl = (Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[519:515]);
  assign Accum2_acc_1895_nl = nl_Accum2_acc_1895_nl[9:0];
  assign nl_Product1_1_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[519:515]));
  assign Product1_1_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1474_nl = ({Accum2_acc_1895_nl , (Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1474_nl = nl_Accum2_acc_1474_nl[15:0];
  assign nl_Accum2_acc_1478_nl = Accum2_acc_1475_nl + Accum2_acc_1474_nl;
  assign Accum2_acc_1478_nl = nl_Accum2_acc_1478_nl[15:0];
  assign nl_Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1479_nl + Accum2_acc_1478_nl;
  assign Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1 = (Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1164:1160]));
  assign Product1_2_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1804:1800]));
  assign Product1_3_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1486_nl = (readslicef_20_16_4(Product1_2_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1486_nl = nl_Accum2_acc_1486_nl[15:0];
  assign nl_Product1_4_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2444:2440]));
  assign Product1_4_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3084:3080]));
  assign Product1_5_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1485_nl = (readslicef_20_16_4(Product1_4_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1485_nl = nl_Accum2_acc_1485_nl[15:0];
  assign nl_Product1_6_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3724:3720]));
  assign Product1_6_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4364:4360]));
  assign Product1_7_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1484_nl = (readslicef_20_16_4(Product1_6_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1484_nl = nl_Accum2_acc_1484_nl[15:0];
  assign nl_Product1_8_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5004:5000]));
  assign Product1_8_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5644:5640]));
  assign Product1_9_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1483_nl = (readslicef_20_16_4(Product1_8_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1483_nl = nl_Accum2_acc_1483_nl[15:0];
  assign nl_Accum2_acc_1492_nl = Accum2_acc_1486_nl + Accum2_acc_1485_nl + Accum2_acc_1484_nl
      + Accum2_acc_1483_nl;
  assign Accum2_acc_1492_nl = nl_Accum2_acc_1492_nl[15:0];
  assign nl_Product1_10_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6284:6280]));
  assign Product1_10_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6924:6920]));
  assign Product1_11_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1482_nl = (readslicef_20_16_4(Product1_10_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1482_nl = nl_Accum2_acc_1482_nl[15:0];
  assign nl_Product1_12_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7564:7560]));
  assign Product1_12_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8204:8200]));
  assign Product1_13_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1481_nl = (readslicef_20_16_4(Product1_12_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1481_nl = nl_Accum2_acc_1481_nl[15:0];
  assign nl_Accum2_acc_1488_nl = Accum2_acc_1482_nl + Accum2_acc_1481_nl;
  assign Accum2_acc_1488_nl = nl_Accum2_acc_1488_nl[15:0];
  assign nl_Accum2_acc_1896_nl = (Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[524:520]);
  assign Accum2_acc_1896_nl = nl_Accum2_acc_1896_nl[9:0];
  assign nl_Product1_1_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[524:520]));
  assign Product1_1_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1487_nl = ({Accum2_acc_1896_nl , (Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1487_nl = nl_Accum2_acc_1487_nl[15:0];
  assign nl_Accum2_acc_1491_nl = Accum2_acc_1488_nl + Accum2_acc_1487_nl;
  assign Accum2_acc_1491_nl = nl_Accum2_acc_1491_nl[15:0];
  assign nl_Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1492_nl + Accum2_acc_1491_nl;
  assign Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1 = (Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1169:1165]));
  assign Product1_2_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1809:1805]));
  assign Product1_3_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1499_nl = (readslicef_20_16_4(Product1_2_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1499_nl = nl_Accum2_acc_1499_nl[15:0];
  assign nl_Product1_4_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2449:2445]));
  assign Product1_4_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3089:3085]));
  assign Product1_5_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1498_nl = (readslicef_20_16_4(Product1_4_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1498_nl = nl_Accum2_acc_1498_nl[15:0];
  assign nl_Product1_6_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3729:3725]));
  assign Product1_6_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4369:4365]));
  assign Product1_7_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1497_nl = (readslicef_20_16_4(Product1_6_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1497_nl = nl_Accum2_acc_1497_nl[15:0];
  assign nl_Product1_8_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5009:5005]));
  assign Product1_8_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5649:5645]));
  assign Product1_9_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1496_nl = (readslicef_20_16_4(Product1_8_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1496_nl = nl_Accum2_acc_1496_nl[15:0];
  assign nl_Accum2_acc_1505_nl = Accum2_acc_1499_nl + Accum2_acc_1498_nl + Accum2_acc_1497_nl
      + Accum2_acc_1496_nl;
  assign Accum2_acc_1505_nl = nl_Accum2_acc_1505_nl[15:0];
  assign nl_Product1_10_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6289:6285]));
  assign Product1_10_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6929:6925]));
  assign Product1_11_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1495_nl = (readslicef_20_16_4(Product1_10_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1495_nl = nl_Accum2_acc_1495_nl[15:0];
  assign nl_Product1_12_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7569:7565]));
  assign Product1_12_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8209:8205]));
  assign Product1_13_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1494_nl = (readslicef_20_16_4(Product1_12_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1494_nl = nl_Accum2_acc_1494_nl[15:0];
  assign nl_Accum2_acc_1501_nl = Accum2_acc_1495_nl + Accum2_acc_1494_nl;
  assign Accum2_acc_1501_nl = nl_Accum2_acc_1501_nl[15:0];
  assign nl_Accum2_acc_1897_nl = (Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[529:525]);
  assign Accum2_acc_1897_nl = nl_Accum2_acc_1897_nl[9:0];
  assign nl_Product1_1_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[529:525]));
  assign Product1_1_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1500_nl = ({Accum2_acc_1897_nl , (Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1500_nl = nl_Accum2_acc_1500_nl[15:0];
  assign nl_Accum2_acc_1504_nl = Accum2_acc_1501_nl + Accum2_acc_1500_nl;
  assign Accum2_acc_1504_nl = nl_Accum2_acc_1504_nl[15:0];
  assign nl_Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1505_nl + Accum2_acc_1504_nl;
  assign Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1 = (Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1174:1170]));
  assign Product1_2_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1814:1810]));
  assign Product1_3_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1512_nl = (readslicef_20_16_4(Product1_2_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1512_nl = nl_Accum2_acc_1512_nl[15:0];
  assign nl_Product1_4_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2454:2450]));
  assign Product1_4_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3094:3090]));
  assign Product1_5_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1511_nl = (readslicef_20_16_4(Product1_4_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1511_nl = nl_Accum2_acc_1511_nl[15:0];
  assign nl_Product1_6_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3734:3730]));
  assign Product1_6_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4374:4370]));
  assign Product1_7_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1510_nl = (readslicef_20_16_4(Product1_6_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1510_nl = nl_Accum2_acc_1510_nl[15:0];
  assign nl_Product1_8_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5014:5010]));
  assign Product1_8_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5654:5650]));
  assign Product1_9_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1509_nl = (readslicef_20_16_4(Product1_8_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1509_nl = nl_Accum2_acc_1509_nl[15:0];
  assign nl_Accum2_acc_1518_nl = Accum2_acc_1512_nl + Accum2_acc_1511_nl + Accum2_acc_1510_nl
      + Accum2_acc_1509_nl;
  assign Accum2_acc_1518_nl = nl_Accum2_acc_1518_nl[15:0];
  assign nl_Product1_10_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6294:6290]));
  assign Product1_10_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6934:6930]));
  assign Product1_11_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1508_nl = (readslicef_20_16_4(Product1_10_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1508_nl = nl_Accum2_acc_1508_nl[15:0];
  assign nl_Product1_12_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7574:7570]));
  assign Product1_12_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8214:8210]));
  assign Product1_13_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1507_nl = (readslicef_20_16_4(Product1_12_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1507_nl = nl_Accum2_acc_1507_nl[15:0];
  assign nl_Accum2_acc_1514_nl = Accum2_acc_1508_nl + Accum2_acc_1507_nl;
  assign Accum2_acc_1514_nl = nl_Accum2_acc_1514_nl[15:0];
  assign nl_Accum2_acc_1898_nl = (Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[534:530]);
  assign Accum2_acc_1898_nl = nl_Accum2_acc_1898_nl[9:0];
  assign nl_Product1_1_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[534:530]));
  assign Product1_1_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1513_nl = ({Accum2_acc_1898_nl , (Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1513_nl = nl_Accum2_acc_1513_nl[15:0];
  assign nl_Accum2_acc_1517_nl = Accum2_acc_1514_nl + Accum2_acc_1513_nl;
  assign Accum2_acc_1517_nl = nl_Accum2_acc_1517_nl[15:0];
  assign nl_Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1518_nl + Accum2_acc_1517_nl;
  assign Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1 = (Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1179:1175]));
  assign Product1_2_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1819:1815]));
  assign Product1_3_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1525_nl = (readslicef_20_16_4(Product1_2_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1525_nl = nl_Accum2_acc_1525_nl[15:0];
  assign nl_Product1_4_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2459:2455]));
  assign Product1_4_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3099:3095]));
  assign Product1_5_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1524_nl = (readslicef_20_16_4(Product1_4_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1524_nl = nl_Accum2_acc_1524_nl[15:0];
  assign nl_Product1_6_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3739:3735]));
  assign Product1_6_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4379:4375]));
  assign Product1_7_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1523_nl = (readslicef_20_16_4(Product1_6_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1523_nl = nl_Accum2_acc_1523_nl[15:0];
  assign nl_Product1_8_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5019:5015]));
  assign Product1_8_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5659:5655]));
  assign Product1_9_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1522_nl = (readslicef_20_16_4(Product1_8_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1522_nl = nl_Accum2_acc_1522_nl[15:0];
  assign nl_Accum2_acc_1531_nl = Accum2_acc_1525_nl + Accum2_acc_1524_nl + Accum2_acc_1523_nl
      + Accum2_acc_1522_nl;
  assign Accum2_acc_1531_nl = nl_Accum2_acc_1531_nl[15:0];
  assign nl_Product1_10_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6299:6295]));
  assign Product1_10_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6939:6935]));
  assign Product1_11_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1521_nl = (readslicef_20_16_4(Product1_10_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1521_nl = nl_Accum2_acc_1521_nl[15:0];
  assign nl_Product1_12_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7579:7575]));
  assign Product1_12_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8219:8215]));
  assign Product1_13_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1520_nl = (readslicef_20_16_4(Product1_12_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1520_nl = nl_Accum2_acc_1520_nl[15:0];
  assign nl_Accum2_acc_1527_nl = Accum2_acc_1521_nl + Accum2_acc_1520_nl;
  assign Accum2_acc_1527_nl = nl_Accum2_acc_1527_nl[15:0];
  assign nl_Accum2_acc_1899_nl = (Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[539:535]);
  assign Accum2_acc_1899_nl = nl_Accum2_acc_1899_nl[9:0];
  assign nl_Product1_1_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[539:535]));
  assign Product1_1_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1526_nl = ({Accum2_acc_1899_nl , (Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1526_nl = nl_Accum2_acc_1526_nl[15:0];
  assign nl_Accum2_acc_1530_nl = Accum2_acc_1527_nl + Accum2_acc_1526_nl;
  assign Accum2_acc_1530_nl = nl_Accum2_acc_1530_nl[15:0];
  assign nl_Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1531_nl + Accum2_acc_1530_nl;
  assign Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1 = (Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1184:1180]));
  assign Product1_2_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1824:1820]));
  assign Product1_3_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1538_nl = (readslicef_20_16_4(Product1_2_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1538_nl = nl_Accum2_acc_1538_nl[15:0];
  assign nl_Product1_4_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2464:2460]));
  assign Product1_4_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3104:3100]));
  assign Product1_5_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1537_nl = (readslicef_20_16_4(Product1_4_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1537_nl = nl_Accum2_acc_1537_nl[15:0];
  assign nl_Product1_6_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3744:3740]));
  assign Product1_6_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4384:4380]));
  assign Product1_7_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1536_nl = (readslicef_20_16_4(Product1_6_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1536_nl = nl_Accum2_acc_1536_nl[15:0];
  assign nl_Product1_8_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5024:5020]));
  assign Product1_8_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5664:5660]));
  assign Product1_9_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1535_nl = (readslicef_20_16_4(Product1_8_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1535_nl = nl_Accum2_acc_1535_nl[15:0];
  assign nl_Accum2_acc_1544_nl = Accum2_acc_1538_nl + Accum2_acc_1537_nl + Accum2_acc_1536_nl
      + Accum2_acc_1535_nl;
  assign Accum2_acc_1544_nl = nl_Accum2_acc_1544_nl[15:0];
  assign nl_Product1_10_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6304:6300]));
  assign Product1_10_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6944:6940]));
  assign Product1_11_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1534_nl = (readslicef_20_16_4(Product1_10_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1534_nl = nl_Accum2_acc_1534_nl[15:0];
  assign nl_Product1_12_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7584:7580]));
  assign Product1_12_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8224:8220]));
  assign Product1_13_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1533_nl = (readslicef_20_16_4(Product1_12_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1533_nl = nl_Accum2_acc_1533_nl[15:0];
  assign nl_Accum2_acc_1540_nl = Accum2_acc_1534_nl + Accum2_acc_1533_nl;
  assign Accum2_acc_1540_nl = nl_Accum2_acc_1540_nl[15:0];
  assign nl_Accum2_acc_1900_nl = (Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[544:540]);
  assign Accum2_acc_1900_nl = nl_Accum2_acc_1900_nl[9:0];
  assign nl_Product1_1_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[544:540]));
  assign Product1_1_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1539_nl = ({Accum2_acc_1900_nl , (Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1539_nl = nl_Accum2_acc_1539_nl[15:0];
  assign nl_Accum2_acc_1543_nl = Accum2_acc_1540_nl + Accum2_acc_1539_nl;
  assign Accum2_acc_1543_nl = nl_Accum2_acc_1543_nl[15:0];
  assign nl_Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1544_nl + Accum2_acc_1543_nl;
  assign Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1 = (Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1189:1185]));
  assign Product1_2_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1829:1825]));
  assign Product1_3_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1551_nl = (readslicef_20_16_4(Product1_2_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1551_nl = nl_Accum2_acc_1551_nl[15:0];
  assign nl_Product1_4_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2469:2465]));
  assign Product1_4_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3109:3105]));
  assign Product1_5_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1550_nl = (readslicef_20_16_4(Product1_4_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1550_nl = nl_Accum2_acc_1550_nl[15:0];
  assign nl_Product1_6_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3749:3745]));
  assign Product1_6_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4389:4385]));
  assign Product1_7_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1549_nl = (readslicef_20_16_4(Product1_6_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1549_nl = nl_Accum2_acc_1549_nl[15:0];
  assign nl_Product1_8_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5029:5025]));
  assign Product1_8_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5669:5665]));
  assign Product1_9_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1548_nl = (readslicef_20_16_4(Product1_8_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1548_nl = nl_Accum2_acc_1548_nl[15:0];
  assign nl_Accum2_acc_1557_nl = Accum2_acc_1551_nl + Accum2_acc_1550_nl + Accum2_acc_1549_nl
      + Accum2_acc_1548_nl;
  assign Accum2_acc_1557_nl = nl_Accum2_acc_1557_nl[15:0];
  assign nl_Product1_10_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6309:6305]));
  assign Product1_10_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6949:6945]));
  assign Product1_11_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1547_nl = (readslicef_20_16_4(Product1_10_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1547_nl = nl_Accum2_acc_1547_nl[15:0];
  assign nl_Product1_12_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7589:7585]));
  assign Product1_12_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8229:8225]));
  assign Product1_13_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1546_nl = (readslicef_20_16_4(Product1_12_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1546_nl = nl_Accum2_acc_1546_nl[15:0];
  assign nl_Accum2_acc_1553_nl = Accum2_acc_1547_nl + Accum2_acc_1546_nl;
  assign Accum2_acc_1553_nl = nl_Accum2_acc_1553_nl[15:0];
  assign nl_Accum2_acc_1901_nl = (Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[549:545]);
  assign Accum2_acc_1901_nl = nl_Accum2_acc_1901_nl[9:0];
  assign nl_Product1_1_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[549:545]));
  assign Product1_1_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1552_nl = ({Accum2_acc_1901_nl , (Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1552_nl = nl_Accum2_acc_1552_nl[15:0];
  assign nl_Accum2_acc_1556_nl = Accum2_acc_1553_nl + Accum2_acc_1552_nl;
  assign Accum2_acc_1556_nl = nl_Accum2_acc_1556_nl[15:0];
  assign nl_Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1557_nl + Accum2_acc_1556_nl;
  assign Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1 = (Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1194:1190]));
  assign Product1_2_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1834:1830]));
  assign Product1_3_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1564_nl = (readslicef_20_16_4(Product1_2_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1564_nl = nl_Accum2_acc_1564_nl[15:0];
  assign nl_Product1_4_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2474:2470]));
  assign Product1_4_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3114:3110]));
  assign Product1_5_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1563_nl = (readslicef_20_16_4(Product1_4_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1563_nl = nl_Accum2_acc_1563_nl[15:0];
  assign nl_Product1_6_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3754:3750]));
  assign Product1_6_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4394:4390]));
  assign Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1562_nl = (readslicef_20_16_4(Product1_6_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1562_nl = nl_Accum2_acc_1562_nl[15:0];
  assign nl_Product1_8_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5034:5030]));
  assign Product1_8_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5674:5670]));
  assign Product1_9_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1561_nl = (readslicef_20_16_4(Product1_8_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1561_nl = nl_Accum2_acc_1561_nl[15:0];
  assign nl_Accum2_acc_1570_nl = Accum2_acc_1564_nl + Accum2_acc_1563_nl + Accum2_acc_1562_nl
      + Accum2_acc_1561_nl;
  assign Accum2_acc_1570_nl = nl_Accum2_acc_1570_nl[15:0];
  assign nl_Product1_10_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6314:6310]));
  assign Product1_10_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6954:6950]));
  assign Product1_11_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1560_nl = (readslicef_20_16_4(Product1_10_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1560_nl = nl_Accum2_acc_1560_nl[15:0];
  assign nl_Product1_12_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7594:7590]));
  assign Product1_12_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8234:8230]));
  assign Product1_13_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1559_nl = (readslicef_20_16_4(Product1_12_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1559_nl = nl_Accum2_acc_1559_nl[15:0];
  assign nl_Accum2_acc_1566_nl = Accum2_acc_1560_nl + Accum2_acc_1559_nl;
  assign Accum2_acc_1566_nl = nl_Accum2_acc_1566_nl[15:0];
  assign nl_Accum2_acc_1902_nl = (Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[554:550]);
  assign Accum2_acc_1902_nl = nl_Accum2_acc_1902_nl[9:0];
  assign nl_Product1_1_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[554:550]));
  assign Product1_1_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1565_nl = ({Accum2_acc_1902_nl , (Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1565_nl = nl_Accum2_acc_1565_nl[15:0];
  assign nl_Accum2_acc_1569_nl = Accum2_acc_1566_nl + Accum2_acc_1565_nl;
  assign Accum2_acc_1569_nl = nl_Accum2_acc_1569_nl[15:0];
  assign nl_Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1570_nl + Accum2_acc_1569_nl;
  assign Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1 = (Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1199:1195]));
  assign Product1_2_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1839:1835]));
  assign Product1_3_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1577_nl = (readslicef_20_16_4(Product1_2_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1577_nl = nl_Accum2_acc_1577_nl[15:0];
  assign nl_Product1_4_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2479:2475]));
  assign Product1_4_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3119:3115]));
  assign Product1_5_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1576_nl = (readslicef_20_16_4(Product1_4_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1576_nl = nl_Accum2_acc_1576_nl[15:0];
  assign nl_Product1_6_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3759:3755]));
  assign Product1_6_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4399:4395]));
  assign Product1_7_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1575_nl = (readslicef_20_16_4(Product1_6_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1575_nl = nl_Accum2_acc_1575_nl[15:0];
  assign nl_Product1_8_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5039:5035]));
  assign Product1_8_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5679:5675]));
  assign Product1_9_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1574_nl = (readslicef_20_16_4(Product1_8_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1574_nl = nl_Accum2_acc_1574_nl[15:0];
  assign nl_Accum2_acc_1583_nl = Accum2_acc_1577_nl + Accum2_acc_1576_nl + Accum2_acc_1575_nl
      + Accum2_acc_1574_nl;
  assign Accum2_acc_1583_nl = nl_Accum2_acc_1583_nl[15:0];
  assign nl_Product1_10_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6319:6315]));
  assign Product1_10_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6959:6955]));
  assign Product1_11_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1573_nl = (readslicef_20_16_4(Product1_10_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1573_nl = nl_Accum2_acc_1573_nl[15:0];
  assign nl_Product1_12_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7599:7595]));
  assign Product1_12_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8239:8235]));
  assign Product1_13_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1572_nl = (readslicef_20_16_4(Product1_12_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1572_nl = nl_Accum2_acc_1572_nl[15:0];
  assign nl_Accum2_acc_1579_nl = Accum2_acc_1573_nl + Accum2_acc_1572_nl;
  assign Accum2_acc_1579_nl = nl_Accum2_acc_1579_nl[15:0];
  assign nl_Accum2_acc_1903_nl = (Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[559:555]);
  assign Accum2_acc_1903_nl = nl_Accum2_acc_1903_nl[9:0];
  assign nl_Product1_1_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[559:555]));
  assign Product1_1_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1578_nl = ({Accum2_acc_1903_nl , (Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1578_nl = nl_Accum2_acc_1578_nl[15:0];
  assign nl_Accum2_acc_1582_nl = Accum2_acc_1579_nl + Accum2_acc_1578_nl;
  assign Accum2_acc_1582_nl = nl_Accum2_acc_1582_nl[15:0];
  assign nl_Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1583_nl + Accum2_acc_1582_nl;
  assign Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1 = (Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1204:1200]));
  assign Product1_2_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1844:1840]));
  assign Product1_3_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1590_nl = (readslicef_20_16_4(Product1_2_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1590_nl = nl_Accum2_acc_1590_nl[15:0];
  assign nl_Product1_4_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2484:2480]));
  assign Product1_4_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3124:3120]));
  assign Product1_5_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1589_nl = (readslicef_20_16_4(Product1_4_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1589_nl = nl_Accum2_acc_1589_nl[15:0];
  assign nl_Product1_6_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3764:3760]));
  assign Product1_6_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4404:4400]));
  assign Product1_7_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1588_nl = (readslicef_20_16_4(Product1_6_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1588_nl = nl_Accum2_acc_1588_nl[15:0];
  assign nl_Product1_8_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5044:5040]));
  assign Product1_8_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5684:5680]));
  assign Product1_9_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1587_nl = (readslicef_20_16_4(Product1_8_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1587_nl = nl_Accum2_acc_1587_nl[15:0];
  assign nl_Accum2_acc_1596_nl = Accum2_acc_1590_nl + Accum2_acc_1589_nl + Accum2_acc_1588_nl
      + Accum2_acc_1587_nl;
  assign Accum2_acc_1596_nl = nl_Accum2_acc_1596_nl[15:0];
  assign nl_Product1_10_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6324:6320]));
  assign Product1_10_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6964:6960]));
  assign Product1_11_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1586_nl = (readslicef_20_16_4(Product1_10_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1586_nl = nl_Accum2_acc_1586_nl[15:0];
  assign nl_Product1_12_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7604:7600]));
  assign Product1_12_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8244:8240]));
  assign Product1_13_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1585_nl = (readslicef_20_16_4(Product1_12_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1585_nl = nl_Accum2_acc_1585_nl[15:0];
  assign nl_Accum2_acc_1592_nl = Accum2_acc_1586_nl + Accum2_acc_1585_nl;
  assign Accum2_acc_1592_nl = nl_Accum2_acc_1592_nl[15:0];
  assign nl_Accum2_acc_1904_nl = (Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[564:560]);
  assign Accum2_acc_1904_nl = nl_Accum2_acc_1904_nl[9:0];
  assign nl_Product1_1_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[564:560]));
  assign Product1_1_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1591_nl = ({Accum2_acc_1904_nl , (Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1591_nl = nl_Accum2_acc_1591_nl[15:0];
  assign nl_Accum2_acc_1595_nl = Accum2_acc_1592_nl + Accum2_acc_1591_nl;
  assign Accum2_acc_1595_nl = nl_Accum2_acc_1595_nl[15:0];
  assign nl_Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1596_nl + Accum2_acc_1595_nl;
  assign Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1 = (Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1209:1205]));
  assign Product1_2_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1849:1845]));
  assign Product1_3_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1603_nl = (readslicef_20_16_4(Product1_2_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1603_nl = nl_Accum2_acc_1603_nl[15:0];
  assign nl_Product1_4_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2489:2485]));
  assign Product1_4_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3129:3125]));
  assign Product1_5_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1602_nl = (readslicef_20_16_4(Product1_4_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1602_nl = nl_Accum2_acc_1602_nl[15:0];
  assign nl_Product1_6_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3769:3765]));
  assign Product1_6_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4409:4405]));
  assign Product1_7_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1601_nl = (readslicef_20_16_4(Product1_6_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1601_nl = nl_Accum2_acc_1601_nl[15:0];
  assign nl_Product1_8_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5049:5045]));
  assign Product1_8_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5689:5685]));
  assign Product1_9_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1600_nl = (readslicef_20_16_4(Product1_8_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1600_nl = nl_Accum2_acc_1600_nl[15:0];
  assign nl_Accum2_acc_1609_nl = Accum2_acc_1603_nl + Accum2_acc_1602_nl + Accum2_acc_1601_nl
      + Accum2_acc_1600_nl;
  assign Accum2_acc_1609_nl = nl_Accum2_acc_1609_nl[15:0];
  assign nl_Product1_10_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6329:6325]));
  assign Product1_10_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6969:6965]));
  assign Product1_11_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1599_nl = (readslicef_20_16_4(Product1_10_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1599_nl = nl_Accum2_acc_1599_nl[15:0];
  assign nl_Product1_12_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7609:7605]));
  assign Product1_12_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8249:8245]));
  assign Product1_13_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1598_nl = (readslicef_20_16_4(Product1_12_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1598_nl = nl_Accum2_acc_1598_nl[15:0];
  assign nl_Accum2_acc_1605_nl = Accum2_acc_1599_nl + Accum2_acc_1598_nl;
  assign Accum2_acc_1605_nl = nl_Accum2_acc_1605_nl[15:0];
  assign nl_Accum2_acc_1905_nl = (Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[569:565]);
  assign Accum2_acc_1905_nl = nl_Accum2_acc_1905_nl[9:0];
  assign nl_Product1_1_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[569:565]));
  assign Product1_1_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1604_nl = ({Accum2_acc_1905_nl , (Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1604_nl = nl_Accum2_acc_1604_nl[15:0];
  assign nl_Accum2_acc_1608_nl = Accum2_acc_1605_nl + Accum2_acc_1604_nl;
  assign Accum2_acc_1608_nl = nl_Accum2_acc_1608_nl[15:0];
  assign nl_Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1609_nl + Accum2_acc_1608_nl;
  assign Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1 = (Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1214:1210]));
  assign Product1_2_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1854:1850]));
  assign Product1_3_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1616_nl = (readslicef_20_16_4(Product1_2_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1616_nl = nl_Accum2_acc_1616_nl[15:0];
  assign nl_Product1_4_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2494:2490]));
  assign Product1_4_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3134:3130]));
  assign Product1_5_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1615_nl = (readslicef_20_16_4(Product1_4_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1615_nl = nl_Accum2_acc_1615_nl[15:0];
  assign nl_Product1_6_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3774:3770]));
  assign Product1_6_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4414:4410]));
  assign Product1_7_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1614_nl = (readslicef_20_16_4(Product1_6_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1614_nl = nl_Accum2_acc_1614_nl[15:0];
  assign nl_Product1_8_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5054:5050]));
  assign Product1_8_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5694:5690]));
  assign Product1_9_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1613_nl = (readslicef_20_16_4(Product1_8_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1613_nl = nl_Accum2_acc_1613_nl[15:0];
  assign nl_Accum2_acc_1622_nl = Accum2_acc_1616_nl + Accum2_acc_1615_nl + Accum2_acc_1614_nl
      + Accum2_acc_1613_nl;
  assign Accum2_acc_1622_nl = nl_Accum2_acc_1622_nl[15:0];
  assign nl_Product1_10_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6334:6330]));
  assign Product1_10_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6974:6970]));
  assign Product1_11_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1612_nl = (readslicef_20_16_4(Product1_10_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1612_nl = nl_Accum2_acc_1612_nl[15:0];
  assign nl_Product1_12_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7614:7610]));
  assign Product1_12_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8254:8250]));
  assign Product1_13_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1611_nl = (readslicef_20_16_4(Product1_12_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1611_nl = nl_Accum2_acc_1611_nl[15:0];
  assign nl_Accum2_acc_1618_nl = Accum2_acc_1612_nl + Accum2_acc_1611_nl;
  assign Accum2_acc_1618_nl = nl_Accum2_acc_1618_nl[15:0];
  assign nl_Accum2_acc_1906_nl = (Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[574:570]);
  assign Accum2_acc_1906_nl = nl_Accum2_acc_1906_nl[9:0];
  assign nl_Product1_1_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[574:570]));
  assign Product1_1_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1617_nl = ({Accum2_acc_1906_nl , (Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1617_nl = nl_Accum2_acc_1617_nl[15:0];
  assign nl_Accum2_acc_1621_nl = Accum2_acc_1618_nl + Accum2_acc_1617_nl;
  assign Accum2_acc_1621_nl = nl_Accum2_acc_1621_nl[15:0];
  assign nl_Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1622_nl + Accum2_acc_1621_nl;
  assign Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1 = (Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1219:1215]));
  assign Product1_2_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1859:1855]));
  assign Product1_3_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1629_nl = (readslicef_20_16_4(Product1_2_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1629_nl = nl_Accum2_acc_1629_nl[15:0];
  assign nl_Product1_4_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2499:2495]));
  assign Product1_4_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3139:3135]));
  assign Product1_5_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1628_nl = (readslicef_20_16_4(Product1_4_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1628_nl = nl_Accum2_acc_1628_nl[15:0];
  assign nl_Product1_6_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3779:3775]));
  assign Product1_6_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4419:4415]));
  assign Product1_7_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1627_nl = (readslicef_20_16_4(Product1_6_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1627_nl = nl_Accum2_acc_1627_nl[15:0];
  assign nl_Product1_8_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5059:5055]));
  assign Product1_8_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5699:5695]));
  assign Product1_9_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1626_nl = (readslicef_20_16_4(Product1_8_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1626_nl = nl_Accum2_acc_1626_nl[15:0];
  assign nl_Accum2_acc_1635_nl = Accum2_acc_1629_nl + Accum2_acc_1628_nl + Accum2_acc_1627_nl
      + Accum2_acc_1626_nl;
  assign Accum2_acc_1635_nl = nl_Accum2_acc_1635_nl[15:0];
  assign nl_Product1_10_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6339:6335]));
  assign Product1_10_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6979:6975]));
  assign Product1_11_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1625_nl = (readslicef_20_16_4(Product1_10_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1625_nl = nl_Accum2_acc_1625_nl[15:0];
  assign nl_Product1_12_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7619:7615]));
  assign Product1_12_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8259:8255]));
  assign Product1_13_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1624_nl = (readslicef_20_16_4(Product1_12_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1624_nl = nl_Accum2_acc_1624_nl[15:0];
  assign nl_Accum2_acc_1631_nl = Accum2_acc_1625_nl + Accum2_acc_1624_nl;
  assign Accum2_acc_1631_nl = nl_Accum2_acc_1631_nl[15:0];
  assign nl_Accum2_acc_1907_nl = (Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[579:575]);
  assign Accum2_acc_1907_nl = nl_Accum2_acc_1907_nl[9:0];
  assign nl_Product1_1_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[579:575]));
  assign Product1_1_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1630_nl = ({Accum2_acc_1907_nl , (Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1630_nl = nl_Accum2_acc_1630_nl[15:0];
  assign nl_Accum2_acc_1634_nl = Accum2_acc_1631_nl + Accum2_acc_1630_nl;
  assign Accum2_acc_1634_nl = nl_Accum2_acc_1634_nl[15:0];
  assign nl_Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1635_nl + Accum2_acc_1634_nl;
  assign Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1 = (Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1224:1220]));
  assign Product1_2_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1864:1860]));
  assign Product1_3_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1642_nl = (readslicef_20_16_4(Product1_2_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1642_nl = nl_Accum2_acc_1642_nl[15:0];
  assign nl_Product1_4_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2504:2500]));
  assign Product1_4_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3144:3140]));
  assign Product1_5_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1641_nl = (readslicef_20_16_4(Product1_4_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1641_nl = nl_Accum2_acc_1641_nl[15:0];
  assign nl_Product1_6_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3784:3780]));
  assign Product1_6_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4424:4420]));
  assign Product1_7_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1640_nl = (readslicef_20_16_4(Product1_6_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1640_nl = nl_Accum2_acc_1640_nl[15:0];
  assign nl_Product1_8_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5064:5060]));
  assign Product1_8_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5704:5700]));
  assign Product1_9_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1639_nl = (readslicef_20_16_4(Product1_8_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1639_nl = nl_Accum2_acc_1639_nl[15:0];
  assign nl_Accum2_acc_1648_nl = Accum2_acc_1642_nl + Accum2_acc_1641_nl + Accum2_acc_1640_nl
      + Accum2_acc_1639_nl;
  assign Accum2_acc_1648_nl = nl_Accum2_acc_1648_nl[15:0];
  assign nl_Product1_10_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6344:6340]));
  assign Product1_10_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6984:6980]));
  assign Product1_11_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1638_nl = (readslicef_20_16_4(Product1_10_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1638_nl = nl_Accum2_acc_1638_nl[15:0];
  assign nl_Product1_12_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7624:7620]));
  assign Product1_12_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8264:8260]));
  assign Product1_13_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1637_nl = (readslicef_20_16_4(Product1_12_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1637_nl = nl_Accum2_acc_1637_nl[15:0];
  assign nl_Accum2_acc_1644_nl = Accum2_acc_1638_nl + Accum2_acc_1637_nl;
  assign Accum2_acc_1644_nl = nl_Accum2_acc_1644_nl[15:0];
  assign nl_Accum2_acc_1908_nl = (Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[584:580]);
  assign Accum2_acc_1908_nl = nl_Accum2_acc_1908_nl[9:0];
  assign nl_Product1_1_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[584:580]));
  assign Product1_1_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1643_nl = ({Accum2_acc_1908_nl , (Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1643_nl = nl_Accum2_acc_1643_nl[15:0];
  assign nl_Accum2_acc_1647_nl = Accum2_acc_1644_nl + Accum2_acc_1643_nl;
  assign Accum2_acc_1647_nl = nl_Accum2_acc_1647_nl[15:0];
  assign nl_Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1648_nl + Accum2_acc_1647_nl;
  assign Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1 = (Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1229:1225]));
  assign Product1_2_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1869:1865]));
  assign Product1_3_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1655_nl = (readslicef_20_16_4(Product1_2_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1655_nl = nl_Accum2_acc_1655_nl[15:0];
  assign nl_Product1_4_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2509:2505]));
  assign Product1_4_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3149:3145]));
  assign Product1_5_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1654_nl = (readslicef_20_16_4(Product1_4_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1654_nl = nl_Accum2_acc_1654_nl[15:0];
  assign nl_Product1_6_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3789:3785]));
  assign Product1_6_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4429:4425]));
  assign Product1_7_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1653_nl = (readslicef_20_16_4(Product1_6_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1653_nl = nl_Accum2_acc_1653_nl[15:0];
  assign nl_Product1_8_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5069:5065]));
  assign Product1_8_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5709:5705]));
  assign Product1_9_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1652_nl = (readslicef_20_16_4(Product1_8_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1652_nl = nl_Accum2_acc_1652_nl[15:0];
  assign nl_Accum2_acc_1661_nl = Accum2_acc_1655_nl + Accum2_acc_1654_nl + Accum2_acc_1653_nl
      + Accum2_acc_1652_nl;
  assign Accum2_acc_1661_nl = nl_Accum2_acc_1661_nl[15:0];
  assign nl_Product1_10_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6349:6345]));
  assign Product1_10_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6989:6985]));
  assign Product1_11_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1651_nl = (readslicef_20_16_4(Product1_10_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1651_nl = nl_Accum2_acc_1651_nl[15:0];
  assign nl_Product1_12_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7629:7625]));
  assign Product1_12_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8269:8265]));
  assign Product1_13_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1650_nl = (readslicef_20_16_4(Product1_12_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1650_nl = nl_Accum2_acc_1650_nl[15:0];
  assign nl_Accum2_acc_1657_nl = Accum2_acc_1651_nl + Accum2_acc_1650_nl;
  assign Accum2_acc_1657_nl = nl_Accum2_acc_1657_nl[15:0];
  assign nl_Accum2_acc_1909_nl = (Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[589:585]);
  assign Accum2_acc_1909_nl = nl_Accum2_acc_1909_nl[9:0];
  assign nl_Product1_1_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[589:585]));
  assign Product1_1_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1656_nl = ({Accum2_acc_1909_nl , (Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1656_nl = nl_Accum2_acc_1656_nl[15:0];
  assign nl_Accum2_acc_1660_nl = Accum2_acc_1657_nl + Accum2_acc_1656_nl;
  assign Accum2_acc_1660_nl = nl_Accum2_acc_1660_nl[15:0];
  assign nl_Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1661_nl + Accum2_acc_1660_nl;
  assign Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1 = (Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1234:1230]));
  assign Product1_2_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1874:1870]));
  assign Product1_3_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1668_nl = (readslicef_20_16_4(Product1_2_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1668_nl = nl_Accum2_acc_1668_nl[15:0];
  assign nl_Product1_4_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2514:2510]));
  assign Product1_4_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3154:3150]));
  assign Product1_5_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1667_nl = (readslicef_20_16_4(Product1_4_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1667_nl = nl_Accum2_acc_1667_nl[15:0];
  assign nl_Product1_6_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3794:3790]));
  assign Product1_6_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4434:4430]));
  assign Product1_7_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1666_nl = (readslicef_20_16_4(Product1_6_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1666_nl = nl_Accum2_acc_1666_nl[15:0];
  assign nl_Product1_8_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5074:5070]));
  assign Product1_8_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5714:5710]));
  assign Product1_9_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1665_nl = (readslicef_20_16_4(Product1_8_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1665_nl = nl_Accum2_acc_1665_nl[15:0];
  assign nl_Accum2_acc_1674_nl = Accum2_acc_1668_nl + Accum2_acc_1667_nl + Accum2_acc_1666_nl
      + Accum2_acc_1665_nl;
  assign Accum2_acc_1674_nl = nl_Accum2_acc_1674_nl[15:0];
  assign nl_Product1_10_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6354:6350]));
  assign Product1_10_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6994:6990]));
  assign Product1_11_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1664_nl = (readslicef_20_16_4(Product1_10_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1664_nl = nl_Accum2_acc_1664_nl[15:0];
  assign nl_Product1_12_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7634:7630]));
  assign Product1_12_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8274:8270]));
  assign Product1_13_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1663_nl = (readslicef_20_16_4(Product1_12_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1663_nl = nl_Accum2_acc_1663_nl[15:0];
  assign nl_Accum2_acc_1670_nl = Accum2_acc_1664_nl + Accum2_acc_1663_nl;
  assign Accum2_acc_1670_nl = nl_Accum2_acc_1670_nl[15:0];
  assign nl_Accum2_acc_1910_nl = (Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[594:590]);
  assign Accum2_acc_1910_nl = nl_Accum2_acc_1910_nl[9:0];
  assign nl_Product1_1_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[594:590]));
  assign Product1_1_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1669_nl = ({Accum2_acc_1910_nl , (Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1669_nl = nl_Accum2_acc_1669_nl[15:0];
  assign nl_Accum2_acc_1673_nl = Accum2_acc_1670_nl + Accum2_acc_1669_nl;
  assign Accum2_acc_1673_nl = nl_Accum2_acc_1673_nl[15:0];
  assign nl_Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1674_nl + Accum2_acc_1673_nl;
  assign Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1 = (Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1239:1235]));
  assign Product1_2_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1879:1875]));
  assign Product1_3_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1681_nl = (readslicef_20_16_4(Product1_2_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1681_nl = nl_Accum2_acc_1681_nl[15:0];
  assign nl_Product1_4_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2519:2515]));
  assign Product1_4_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3159:3155]));
  assign Product1_5_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1680_nl = (readslicef_20_16_4(Product1_4_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1680_nl = nl_Accum2_acc_1680_nl[15:0];
  assign nl_Product1_6_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3799:3795]));
  assign Product1_6_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4439:4435]));
  assign Product1_7_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1679_nl = (readslicef_20_16_4(Product1_6_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1679_nl = nl_Accum2_acc_1679_nl[15:0];
  assign nl_Product1_8_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5079:5075]));
  assign Product1_8_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5719:5715]));
  assign Product1_9_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1678_nl = (readslicef_20_16_4(Product1_8_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1678_nl = nl_Accum2_acc_1678_nl[15:0];
  assign nl_Accum2_acc_1687_nl = Accum2_acc_1681_nl + Accum2_acc_1680_nl + Accum2_acc_1679_nl
      + Accum2_acc_1678_nl;
  assign Accum2_acc_1687_nl = nl_Accum2_acc_1687_nl[15:0];
  assign nl_Product1_10_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6359:6355]));
  assign Product1_10_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[6999:6995]));
  assign Product1_11_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1677_nl = (readslicef_20_16_4(Product1_10_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1677_nl = nl_Accum2_acc_1677_nl[15:0];
  assign nl_Product1_12_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7639:7635]));
  assign Product1_12_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8279:8275]));
  assign Product1_13_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1676_nl = (readslicef_20_16_4(Product1_12_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1676_nl = nl_Accum2_acc_1676_nl[15:0];
  assign nl_Accum2_acc_1683_nl = Accum2_acc_1677_nl + Accum2_acc_1676_nl;
  assign Accum2_acc_1683_nl = nl_Accum2_acc_1683_nl[15:0];
  assign nl_Accum2_acc_1911_nl = (Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[599:595]);
  assign Accum2_acc_1911_nl = nl_Accum2_acc_1911_nl[9:0];
  assign nl_Product1_1_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[599:595]));
  assign Product1_1_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1682_nl = ({Accum2_acc_1911_nl , (Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1682_nl = nl_Accum2_acc_1682_nl[15:0];
  assign nl_Accum2_acc_1686_nl = Accum2_acc_1683_nl + Accum2_acc_1682_nl;
  assign Accum2_acc_1686_nl = nl_Accum2_acc_1686_nl[15:0];
  assign nl_Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1687_nl + Accum2_acc_1686_nl;
  assign Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1 = (Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1244:1240]));
  assign Product1_2_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1884:1880]));
  assign Product1_3_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1694_nl = (readslicef_20_16_4(Product1_2_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1694_nl = nl_Accum2_acc_1694_nl[15:0];
  assign nl_Product1_4_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2524:2520]));
  assign Product1_4_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3164:3160]));
  assign Product1_5_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1693_nl = (readslicef_20_16_4(Product1_4_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1693_nl = nl_Accum2_acc_1693_nl[15:0];
  assign nl_Product1_6_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3804:3800]));
  assign Product1_6_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4444:4440]));
  assign Product1_7_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1692_nl = (readslicef_20_16_4(Product1_6_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1692_nl = nl_Accum2_acc_1692_nl[15:0];
  assign nl_Product1_8_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5084:5080]));
  assign Product1_8_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5724:5720]));
  assign Product1_9_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1691_nl = (readslicef_20_16_4(Product1_8_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1691_nl = nl_Accum2_acc_1691_nl[15:0];
  assign nl_Accum2_acc_1700_nl = Accum2_acc_1694_nl + Accum2_acc_1693_nl + Accum2_acc_1692_nl
      + Accum2_acc_1691_nl;
  assign Accum2_acc_1700_nl = nl_Accum2_acc_1700_nl[15:0];
  assign nl_Product1_10_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6364:6360]));
  assign Product1_10_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7004:7000]));
  assign Product1_11_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1690_nl = (readslicef_20_16_4(Product1_10_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1690_nl = nl_Accum2_acc_1690_nl[15:0];
  assign nl_Product1_12_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7644:7640]));
  assign Product1_12_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8284:8280]));
  assign Product1_13_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1689_nl = (readslicef_20_16_4(Product1_12_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1689_nl = nl_Accum2_acc_1689_nl[15:0];
  assign nl_Accum2_acc_1696_nl = Accum2_acc_1690_nl + Accum2_acc_1689_nl;
  assign Accum2_acc_1696_nl = nl_Accum2_acc_1696_nl[15:0];
  assign nl_Accum2_acc_1912_nl = (Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[604:600]);
  assign Accum2_acc_1912_nl = nl_Accum2_acc_1912_nl[9:0];
  assign nl_Product1_1_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[604:600]));
  assign Product1_1_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1695_nl = ({Accum2_acc_1912_nl , (Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1695_nl = nl_Accum2_acc_1695_nl[15:0];
  assign nl_Accum2_acc_1699_nl = Accum2_acc_1696_nl + Accum2_acc_1695_nl;
  assign Accum2_acc_1699_nl = nl_Accum2_acc_1699_nl[15:0];
  assign nl_Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1700_nl + Accum2_acc_1699_nl;
  assign Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1 = (Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1249:1245]));
  assign Product1_2_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1889:1885]));
  assign Product1_3_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1707_nl = (readslicef_20_16_4(Product1_2_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1707_nl = nl_Accum2_acc_1707_nl[15:0];
  assign nl_Product1_4_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2529:2525]));
  assign Product1_4_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3169:3165]));
  assign Product1_5_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1706_nl = (readslicef_20_16_4(Product1_4_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1706_nl = nl_Accum2_acc_1706_nl[15:0];
  assign nl_Product1_6_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3809:3805]));
  assign Product1_6_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4449:4445]));
  assign Product1_7_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1705_nl = (readslicef_20_16_4(Product1_6_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1705_nl = nl_Accum2_acc_1705_nl[15:0];
  assign nl_Product1_8_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5089:5085]));
  assign Product1_8_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5729:5725]));
  assign Product1_9_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1704_nl = (readslicef_20_16_4(Product1_8_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1704_nl = nl_Accum2_acc_1704_nl[15:0];
  assign nl_Accum2_acc_1713_nl = Accum2_acc_1707_nl + Accum2_acc_1706_nl + Accum2_acc_1705_nl
      + Accum2_acc_1704_nl;
  assign Accum2_acc_1713_nl = nl_Accum2_acc_1713_nl[15:0];
  assign nl_Product1_10_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6369:6365]));
  assign Product1_10_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7009:7005]));
  assign Product1_11_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1703_nl = (readslicef_20_16_4(Product1_10_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1703_nl = nl_Accum2_acc_1703_nl[15:0];
  assign nl_Product1_12_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7649:7645]));
  assign Product1_12_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8289:8285]));
  assign Product1_13_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1702_nl = (readslicef_20_16_4(Product1_12_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1702_nl = nl_Accum2_acc_1702_nl[15:0];
  assign nl_Accum2_acc_1709_nl = Accum2_acc_1703_nl + Accum2_acc_1702_nl;
  assign Accum2_acc_1709_nl = nl_Accum2_acc_1709_nl[15:0];
  assign nl_Accum2_acc_1913_nl = (Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[609:605]);
  assign Accum2_acc_1913_nl = nl_Accum2_acc_1913_nl[9:0];
  assign nl_Product1_1_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[609:605]));
  assign Product1_1_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1708_nl = ({Accum2_acc_1913_nl , (Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1708_nl = nl_Accum2_acc_1708_nl[15:0];
  assign nl_Accum2_acc_1712_nl = Accum2_acc_1709_nl + Accum2_acc_1708_nl;
  assign Accum2_acc_1712_nl = nl_Accum2_acc_1712_nl[15:0];
  assign nl_Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1713_nl + Accum2_acc_1712_nl;
  assign Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1 = (Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1254:1250]));
  assign Product1_2_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1894:1890]));
  assign Product1_3_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1720_nl = (readslicef_20_16_4(Product1_2_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1720_nl = nl_Accum2_acc_1720_nl[15:0];
  assign nl_Product1_4_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2534:2530]));
  assign Product1_4_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3174:3170]));
  assign Product1_5_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1719_nl = (readslicef_20_16_4(Product1_4_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1719_nl = nl_Accum2_acc_1719_nl[15:0];
  assign nl_Product1_6_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3814:3810]));
  assign Product1_6_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4454:4450]));
  assign Product1_7_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1718_nl = (readslicef_20_16_4(Product1_6_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1718_nl = nl_Accum2_acc_1718_nl[15:0];
  assign nl_Product1_8_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5094:5090]));
  assign Product1_8_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5734:5730]));
  assign Product1_9_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1717_nl = (readslicef_20_16_4(Product1_8_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1717_nl = nl_Accum2_acc_1717_nl[15:0];
  assign nl_Accum2_acc_1726_nl = Accum2_acc_1720_nl + Accum2_acc_1719_nl + Accum2_acc_1718_nl
      + Accum2_acc_1717_nl;
  assign Accum2_acc_1726_nl = nl_Accum2_acc_1726_nl[15:0];
  assign nl_Product1_10_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6374:6370]));
  assign Product1_10_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7014:7010]));
  assign Product1_11_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1716_nl = (readslicef_20_16_4(Product1_10_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1716_nl = nl_Accum2_acc_1716_nl[15:0];
  assign nl_Product1_12_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7654:7650]));
  assign Product1_12_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8294:8290]));
  assign Product1_13_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1715_nl = (readslicef_20_16_4(Product1_12_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1715_nl = nl_Accum2_acc_1715_nl[15:0];
  assign nl_Accum2_acc_1722_nl = Accum2_acc_1716_nl + Accum2_acc_1715_nl;
  assign Accum2_acc_1722_nl = nl_Accum2_acc_1722_nl[15:0];
  assign nl_Accum2_acc_1914_nl = (Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[614:610]);
  assign Accum2_acc_1914_nl = nl_Accum2_acc_1914_nl[9:0];
  assign nl_Product1_1_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[614:610]));
  assign Product1_1_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1721_nl = ({Accum2_acc_1914_nl , (Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1721_nl = nl_Accum2_acc_1721_nl[15:0];
  assign nl_Accum2_acc_1725_nl = Accum2_acc_1722_nl + Accum2_acc_1721_nl;
  assign Accum2_acc_1725_nl = nl_Accum2_acc_1725_nl[15:0];
  assign nl_Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1726_nl + Accum2_acc_1725_nl;
  assign Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1 = (Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1259:1255]));
  assign Product1_2_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1899:1895]));
  assign Product1_3_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1733_nl = (readslicef_20_16_4(Product1_2_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1733_nl = nl_Accum2_acc_1733_nl[15:0];
  assign nl_Product1_4_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2539:2535]));
  assign Product1_4_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3179:3175]));
  assign Product1_5_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1732_nl = (readslicef_20_16_4(Product1_4_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1732_nl = nl_Accum2_acc_1732_nl[15:0];
  assign nl_Product1_6_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3819:3815]));
  assign Product1_6_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4459:4455]));
  assign Product1_7_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1731_nl = (readslicef_20_16_4(Product1_6_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1731_nl = nl_Accum2_acc_1731_nl[15:0];
  assign nl_Product1_8_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5099:5095]));
  assign Product1_8_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5739:5735]));
  assign Product1_9_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1730_nl = (readslicef_20_16_4(Product1_8_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1730_nl = nl_Accum2_acc_1730_nl[15:0];
  assign nl_Accum2_acc_1739_nl = Accum2_acc_1733_nl + Accum2_acc_1732_nl + Accum2_acc_1731_nl
      + Accum2_acc_1730_nl;
  assign Accum2_acc_1739_nl = nl_Accum2_acc_1739_nl[15:0];
  assign nl_Product1_10_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6379:6375]));
  assign Product1_10_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7019:7015]));
  assign Product1_11_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1729_nl = (readslicef_20_16_4(Product1_10_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1729_nl = nl_Accum2_acc_1729_nl[15:0];
  assign nl_Product1_12_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7659:7655]));
  assign Product1_12_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8299:8295]));
  assign Product1_13_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1728_nl = (readslicef_20_16_4(Product1_12_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1728_nl = nl_Accum2_acc_1728_nl[15:0];
  assign nl_Accum2_acc_1735_nl = Accum2_acc_1729_nl + Accum2_acc_1728_nl;
  assign Accum2_acc_1735_nl = nl_Accum2_acc_1735_nl[15:0];
  assign nl_Accum2_acc_1915_nl = (Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[619:615]);
  assign Accum2_acc_1915_nl = nl_Accum2_acc_1915_nl[9:0];
  assign nl_Product1_1_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[619:615]));
  assign Product1_1_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1734_nl = ({Accum2_acc_1915_nl , (Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1734_nl = nl_Accum2_acc_1734_nl[15:0];
  assign nl_Accum2_acc_1738_nl = Accum2_acc_1735_nl + Accum2_acc_1734_nl;
  assign Accum2_acc_1738_nl = nl_Accum2_acc_1738_nl[15:0];
  assign nl_Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1739_nl + Accum2_acc_1738_nl;
  assign Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1 = (Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1264:1260]));
  assign Product1_2_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1904:1900]));
  assign Product1_3_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1746_nl = (readslicef_20_16_4(Product1_2_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1746_nl = nl_Accum2_acc_1746_nl[15:0];
  assign nl_Product1_4_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2544:2540]));
  assign Product1_4_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3184:3180]));
  assign Product1_5_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1745_nl = (readslicef_20_16_4(Product1_4_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1745_nl = nl_Accum2_acc_1745_nl[15:0];
  assign nl_Product1_6_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3824:3820]));
  assign Product1_6_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4464:4460]));
  assign Product1_7_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1744_nl = (readslicef_20_16_4(Product1_6_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1744_nl = nl_Accum2_acc_1744_nl[15:0];
  assign nl_Product1_8_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5104:5100]));
  assign Product1_8_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5744:5740]));
  assign Product1_9_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1743_nl = (readslicef_20_16_4(Product1_8_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1743_nl = nl_Accum2_acc_1743_nl[15:0];
  assign nl_Accum2_acc_1752_nl = Accum2_acc_1746_nl + Accum2_acc_1745_nl + Accum2_acc_1744_nl
      + Accum2_acc_1743_nl;
  assign Accum2_acc_1752_nl = nl_Accum2_acc_1752_nl[15:0];
  assign nl_Product1_10_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6384:6380]));
  assign Product1_10_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7024:7020]));
  assign Product1_11_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1742_nl = (readslicef_20_16_4(Product1_10_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1742_nl = nl_Accum2_acc_1742_nl[15:0];
  assign nl_Product1_12_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7664:7660]));
  assign Product1_12_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8304:8300]));
  assign Product1_13_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1741_nl = (readslicef_20_16_4(Product1_12_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1741_nl = nl_Accum2_acc_1741_nl[15:0];
  assign nl_Accum2_acc_1748_nl = Accum2_acc_1742_nl + Accum2_acc_1741_nl;
  assign Accum2_acc_1748_nl = nl_Accum2_acc_1748_nl[15:0];
  assign nl_Accum2_acc_1916_nl = (Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[624:620]);
  assign Accum2_acc_1916_nl = nl_Accum2_acc_1916_nl[9:0];
  assign nl_Product1_1_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[624:620]));
  assign Product1_1_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1747_nl = ({Accum2_acc_1916_nl , (Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1747_nl = nl_Accum2_acc_1747_nl[15:0];
  assign nl_Accum2_acc_1751_nl = Accum2_acc_1748_nl + Accum2_acc_1747_nl;
  assign Accum2_acc_1751_nl = nl_Accum2_acc_1751_nl[15:0];
  assign nl_Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1752_nl + Accum2_acc_1751_nl;
  assign Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1 = (Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1269:1265]));
  assign Product1_2_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1909:1905]));
  assign Product1_3_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1759_nl = (readslicef_20_16_4(Product1_2_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1759_nl = nl_Accum2_acc_1759_nl[15:0];
  assign nl_Product1_4_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2549:2545]));
  assign Product1_4_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3189:3185]));
  assign Product1_5_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1758_nl = (readslicef_20_16_4(Product1_4_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1758_nl = nl_Accum2_acc_1758_nl[15:0];
  assign nl_Product1_6_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3829:3825]));
  assign Product1_6_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4469:4465]));
  assign Product1_7_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1757_nl = (readslicef_20_16_4(Product1_6_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1757_nl = nl_Accum2_acc_1757_nl[15:0];
  assign nl_Product1_8_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5109:5105]));
  assign Product1_8_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5749:5745]));
  assign Product1_9_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1756_nl = (readslicef_20_16_4(Product1_8_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1756_nl = nl_Accum2_acc_1756_nl[15:0];
  assign nl_Accum2_acc_1765_nl = Accum2_acc_1759_nl + Accum2_acc_1758_nl + Accum2_acc_1757_nl
      + Accum2_acc_1756_nl;
  assign Accum2_acc_1765_nl = nl_Accum2_acc_1765_nl[15:0];
  assign nl_Product1_10_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6389:6385]));
  assign Product1_10_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7029:7025]));
  assign Product1_11_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1755_nl = (readslicef_20_16_4(Product1_10_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1755_nl = nl_Accum2_acc_1755_nl[15:0];
  assign nl_Product1_12_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7669:7665]));
  assign Product1_12_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8309:8305]));
  assign Product1_13_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1754_nl = (readslicef_20_16_4(Product1_12_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1754_nl = nl_Accum2_acc_1754_nl[15:0];
  assign nl_Accum2_acc_1761_nl = Accum2_acc_1755_nl + Accum2_acc_1754_nl;
  assign Accum2_acc_1761_nl = nl_Accum2_acc_1761_nl[15:0];
  assign nl_Accum2_acc_1917_nl = (Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[629:625]);
  assign Accum2_acc_1917_nl = nl_Accum2_acc_1917_nl[9:0];
  assign nl_Product1_1_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[629:625]));
  assign Product1_1_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1760_nl = ({Accum2_acc_1917_nl , (Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1760_nl = nl_Accum2_acc_1760_nl[15:0];
  assign nl_Accum2_acc_1764_nl = Accum2_acc_1761_nl + Accum2_acc_1760_nl;
  assign Accum2_acc_1764_nl = nl_Accum2_acc_1764_nl[15:0];
  assign nl_Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1765_nl + Accum2_acc_1764_nl;
  assign Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1 = (Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1274:1270]));
  assign Product1_2_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1914:1910]));
  assign Product1_3_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1772_nl = (readslicef_20_16_4(Product1_2_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1772_nl = nl_Accum2_acc_1772_nl[15:0];
  assign nl_Product1_4_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2554:2550]));
  assign Product1_4_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3194:3190]));
  assign Product1_5_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1771_nl = (readslicef_20_16_4(Product1_4_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1771_nl = nl_Accum2_acc_1771_nl[15:0];
  assign nl_Product1_6_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3834:3830]));
  assign Product1_6_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4474:4470]));
  assign Product1_7_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1770_nl = (readslicef_20_16_4(Product1_6_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1770_nl = nl_Accum2_acc_1770_nl[15:0];
  assign nl_Product1_8_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5114:5110]));
  assign Product1_8_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5754:5750]));
  assign Product1_9_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1769_nl = (readslicef_20_16_4(Product1_8_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1769_nl = nl_Accum2_acc_1769_nl[15:0];
  assign nl_Accum2_acc_1778_nl = Accum2_acc_1772_nl + Accum2_acc_1771_nl + Accum2_acc_1770_nl
      + Accum2_acc_1769_nl;
  assign Accum2_acc_1778_nl = nl_Accum2_acc_1778_nl[15:0];
  assign nl_Product1_10_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6394:6390]));
  assign Product1_10_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7034:7030]));
  assign Product1_11_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1768_nl = (readslicef_20_16_4(Product1_10_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1768_nl = nl_Accum2_acc_1768_nl[15:0];
  assign nl_Product1_12_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7674:7670]));
  assign Product1_12_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8314:8310]));
  assign Product1_13_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1767_nl = (readslicef_20_16_4(Product1_12_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1767_nl = nl_Accum2_acc_1767_nl[15:0];
  assign nl_Accum2_acc_1774_nl = Accum2_acc_1768_nl + Accum2_acc_1767_nl;
  assign Accum2_acc_1774_nl = nl_Accum2_acc_1774_nl[15:0];
  assign nl_Accum2_acc_1918_nl = (Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[634:630]);
  assign Accum2_acc_1918_nl = nl_Accum2_acc_1918_nl[9:0];
  assign nl_Product1_1_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[634:630]));
  assign Product1_1_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1773_nl = ({Accum2_acc_1918_nl , (Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1773_nl = nl_Accum2_acc_1773_nl[15:0];
  assign nl_Accum2_acc_1777_nl = Accum2_acc_1774_nl + Accum2_acc_1773_nl;
  assign Accum2_acc_1777_nl = nl_Accum2_acc_1777_nl[15:0];
  assign nl_Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1778_nl + Accum2_acc_1777_nl;
  assign Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 = (Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[14:10]!=5'b00000);
  assign nl_Product1_2_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[31:16])) * $signed((w2_rsci_idat[1279:1275]));
  assign Product1_2_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_2_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_3_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[47:32])) * $signed((w2_rsci_idat[1919:1915]));
  assign Product1_3_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_3_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1785_nl = (readslicef_20_16_4(Product1_2_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_3_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1785_nl = nl_Accum2_acc_1785_nl[15:0];
  assign nl_Product1_4_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[63:48])) * $signed((w2_rsci_idat[2559:2555]));
  assign Product1_4_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_4_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_5_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[79:64])) * $signed((w2_rsci_idat[3199:3195]));
  assign Product1_5_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_5_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1784_nl = (readslicef_20_16_4(Product1_4_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_5_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1784_nl = nl_Accum2_acc_1784_nl[15:0];
  assign nl_Product1_6_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[95:80])) * $signed((w2_rsci_idat[3839:3835]));
  assign Product1_6_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_6_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_7_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[111:96])) * $signed((w2_rsci_idat[4479:4475]));
  assign Product1_7_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_7_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1783_nl = (readslicef_20_16_4(Product1_6_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_7_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1783_nl = nl_Accum2_acc_1783_nl[15:0];
  assign nl_Product1_8_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[127:112])) * $signed((w2_rsci_idat[5119:5115]));
  assign Product1_8_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_8_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_9_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[143:128])) * $signed((w2_rsci_idat[5759:5755]));
  assign Product1_9_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_9_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1782_nl = (readslicef_20_16_4(Product1_8_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_9_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1782_nl = nl_Accum2_acc_1782_nl[15:0];
  assign nl_Accum2_acc_1791_nl = Accum2_acc_1785_nl + Accum2_acc_1784_nl + Accum2_acc_1783_nl
      + Accum2_acc_1782_nl;
  assign Accum2_acc_1791_nl = nl_Accum2_acc_1791_nl[15:0];
  assign nl_Product1_10_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[159:144])) * $signed((w2_rsci_idat[6399:6395]));
  assign Product1_10_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_10_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_11_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[175:160])) * $signed((w2_rsci_idat[7039:7035]));
  assign Product1_11_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_11_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1781_nl = (readslicef_20_16_4(Product1_10_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_11_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1781_nl = nl_Accum2_acc_1781_nl[15:0];
  assign nl_Product1_12_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[191:176])) * $signed((w2_rsci_idat[7679:7675]));
  assign Product1_12_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_12_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Product1_13_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[207:192])) * $signed((w2_rsci_idat[8319:8315]));
  assign Product1_13_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_13_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1780_nl = (readslicef_20_16_4(Product1_12_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl))
      + (readslicef_20_16_4(Product1_13_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1780_nl = nl_Accum2_acc_1780_nl[15:0];
  assign nl_Accum2_acc_1787_nl = Accum2_acc_1781_nl + Accum2_acc_1780_nl;
  assign Accum2_acc_1787_nl = nl_Accum2_acc_1787_nl[15:0];
  assign nl_Accum2_acc_1919_nl = (Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[639:635]);
  assign Accum2_acc_1919_nl = nl_Accum2_acc_1919_nl[9:0];
  assign nl_Product1_1_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[15:0])) * $signed((w2_rsci_idat[639:635]));
  assign Product1_1_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_1_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign nl_Accum2_acc_1786_nl = ({Accum2_acc_1919_nl , (Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(Product1_1_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl));
  assign Accum2_acc_1786_nl = nl_Accum2_acc_1786_nl[15:0];
  assign nl_Accum2_acc_1790_nl = Accum2_acc_1787_nl + Accum2_acc_1786_nl;
  assign Accum2_acc_1790_nl = nl_Accum2_acc_1790_nl[15:0];
  assign nl_Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1 = Accum2_acc_1791_nl + Accum2_acc_1790_nl;
  assign Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1 = nl_Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[15:0];
  assign nl_Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_0}))
      * $signed((w5_rsci_idat[1604:1600]));
  assign Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1
      = readslicef_15_11_4(Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl);
  assign nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_193_9 , layer4_out_conc_193_8_1 ,
      layer4_out_conc_193_0})) * $signed((w5_rsci_idat[4:0]));
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1
      = readslicef_15_11_4(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl);
  assign nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_193_9 , layer4_out_conc_193_8_1 ,
      layer4_out_conc_193_0})) * $signed((w5_rsci_idat[9:5]));
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1
      = readslicef_15_11_4(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl
      =  -conv_s2s_16_17(nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nl_Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8959:8955]));
  assign Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_128_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8954:8950]));
  assign Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_127_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8949:8945]));
  assign Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_126_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8944:8940]));
  assign Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_125_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8939:8935]));
  assign Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_124_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8934:8930]));
  assign Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_123_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8929:8925]));
  assign Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_122_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8924:8920]));
  assign Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_121_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8919:8915]));
  assign Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_120_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8914:8910]));
  assign Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_119_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8909:8905]));
  assign Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_118_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8904:8900]));
  assign Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_117_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8899:8895]));
  assign Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_116_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8894:8890]));
  assign Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_115_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8889:8885]));
  assign Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_114_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8884:8880]));
  assign Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_113_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8879:8875]));
  assign Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_112_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8874:8870]));
  assign Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_111_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8869:8865]));
  assign Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_110_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8864:8860]));
  assign Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_109_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8859:8855]));
  assign Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_108_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8854:8850]));
  assign Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_107_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8849:8845]));
  assign Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_106_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8844:8840]));
  assign Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_105_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8839:8835]));
  assign Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_104_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8834:8830]));
  assign Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_103_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8829:8825]));
  assign Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_102_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8824:8820]));
  assign Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_101_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8819:8815]));
  assign Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_100_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8814:8810]));
  assign Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_99_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8809:8805]));
  assign Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_98_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8804:8800]));
  assign Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_97_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8799:8795]));
  assign Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_96_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8794:8790]));
  assign Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_95_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8789:8785]));
  assign Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_94_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8784:8780]));
  assign Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_93_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8779:8775]));
  assign Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_92_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8774:8770]));
  assign Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_91_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8769:8765]));
  assign Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_90_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8764:8760]));
  assign Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_89_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8759:8755]));
  assign Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_88_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8754:8750]));
  assign Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_87_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8749:8745]));
  assign Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_86_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8744:8740]));
  assign Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_85_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8739:8735]));
  assign Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_84_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8734:8730]));
  assign Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_83_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8729:8725]));
  assign Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_82_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8724:8720]));
  assign Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_81_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8719:8715]));
  assign Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_80_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8714:8710]));
  assign Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_79_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8709:8705]));
  assign Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_78_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8704:8700]));
  assign Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_77_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8699:8695]));
  assign Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_76_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8694:8690]));
  assign Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_75_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8689:8685]));
  assign Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_74_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8684:8680]));
  assign Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_73_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8679:8675]));
  assign Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_72_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8674:8670]));
  assign Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_71_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8669:8665]));
  assign Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_70_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8664:8660]));
  assign Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_69_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8659:8655]));
  assign Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_68_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8654:8650]));
  assign Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_67_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8649:8645]));
  assign Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_66_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8644:8640]));
  assign Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_65_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8639:8635]));
  assign Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_64_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8634:8630]));
  assign Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_63_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8629:8625]));
  assign Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_62_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8624:8620]));
  assign Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_61_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8619:8615]));
  assign Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_60_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8614:8610]));
  assign Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_59_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8609:8605]));
  assign Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_58_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8604:8600]));
  assign Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_57_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8599:8595]));
  assign Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_56_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8594:8590]));
  assign Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_55_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8589:8585]));
  assign Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_54_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8584:8580]));
  assign Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_53_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8579:8575]));
  assign Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_52_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8574:8570]));
  assign Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_51_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8569:8565]));
  assign Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_50_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8564:8560]));
  assign Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_49_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8559:8555]));
  assign Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_48_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8554:8550]));
  assign Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_47_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8549:8545]));
  assign Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_46_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8544:8540]));
  assign Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_45_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8539:8535]));
  assign Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_44_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8534:8530]));
  assign Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_43_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8529:8525]));
  assign Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_42_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8524:8520]));
  assign Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_41_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8519:8515]));
  assign Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_40_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8514:8510]));
  assign Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_39_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8509:8505]));
  assign Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_38_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8504:8500]));
  assign Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_37_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8499:8495]));
  assign Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_36_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8494:8490]));
  assign Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_35_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8489:8485]));
  assign Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_34_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8484:8480]));
  assign Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_33_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8479:8475]));
  assign Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_32_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8474:8470]));
  assign Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_31_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8469:8465]));
  assign Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_30_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8464:8460]));
  assign Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_29_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8459:8455]));
  assign Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_28_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8454:8450]));
  assign Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_27_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8449:8445]));
  assign Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_26_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8444:8440]));
  assign Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_25_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8439:8435]));
  assign Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_24_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8434:8430]));
  assign Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_23_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8429:8425]));
  assign Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_22_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8424:8420]));
  assign Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_21_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8419:8415]));
  assign Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_20_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8414:8410]));
  assign Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_19_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8409:8405]));
  assign Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_18_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8404:8400]));
  assign Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_17_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8399:8395]));
  assign Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_16_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8394:8390]));
  assign Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_15_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8389:8385]));
  assign Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_14_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8384:8380]));
  assign Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_13_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8379:8375]));
  assign Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_12_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8374:8370]));
  assign Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_11_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8369:8365]));
  assign Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_10_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8364:8360]));
  assign Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_9_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8359:8355]));
  assign Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_8_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8354:8350]));
  assign Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_7_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8349:8345]));
  assign Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_6_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8344:8340]));
  assign Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_5_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8339:8335]));
  assign Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_4_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8334:8330]));
  assign Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_3_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8329:8325]));
  assign Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_2_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nl_Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = $signed((input_1_rsci_idat[223:208])) * $signed((w2_rsci_idat[8324:8320]));
  assign Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl
      = nl_Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl[19:0];
  assign Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_itm_19_4_1
      = readslicef_20_16_4(Product1_14_Product2_1_nnet_product_mult_input_t_config2_weight_t_product_mul_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9 = ((Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_0 = ((Accum1_14_Accum2_105_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9 = ((Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_0 = ((Accum1_14_Accum2_106_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9 = ((Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_0 = ((Accum1_14_Accum2_126_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9 = ((Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_0 = ((Accum1_14_Accum2_127_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9 = ((Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_0 = ((Accum1_14_Accum2_128_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9 = ((Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_0 = ((Accum1_14_Accum2_124_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9 = ((Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_0 = ((Accum1_14_Accum2_125_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9 = ((Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_0 = ((Accum1_14_Accum2_122_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9 = ((Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_0 = ((Accum1_14_Accum2_123_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9 = ((Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_0 = ((Accum1_14_Accum2_120_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9 = ((Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_0 = ((Accum1_14_Accum2_121_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9 = ((Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_0 = ((Accum1_14_Accum2_118_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9 = ((Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_0 = ((Accum1_14_Accum2_119_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9 = ((Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_0 = ((Accum1_14_Accum2_116_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9 = ((Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_0 = ((Accum1_14_Accum2_117_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9 = ((Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_0 = ((Accum1_14_Accum2_114_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9 = ((Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_0 = ((Accum1_14_Accum2_115_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9 = ((Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_0 = ((Accum1_14_Accum2_112_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9 = ((Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_0 = ((Accum1_14_Accum2_113_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9 = ((Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_0 = ((Accum1_14_Accum2_110_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9 = ((Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_0 = ((Accum1_14_Accum2_111_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9 = ((Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_0 = ((Accum1_14_Accum2_108_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9 = ((Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_0 = ((Accum1_14_Accum2_109_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_193_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1);
  assign layer4_out_conc_193_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_193_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_0_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_195_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1);
  assign layer4_out_conc_195_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_195_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_1_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_197_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1);
  assign layer4_out_conc_197_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_197_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_2_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_199_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1);
  assign layer4_out_conc_199_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_199_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_3_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_201_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1);
  assign layer4_out_conc_201_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_201_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_4_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_203_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1);
  assign layer4_out_conc_203_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_203_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_5_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_205_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1);
  assign layer4_out_conc_205_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_205_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_6_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_207_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1);
  assign layer4_out_conc_207_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_207_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_7_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_209_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1);
  assign layer4_out_conc_209_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_209_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_8_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_211_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1);
  assign layer4_out_conc_211_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_211_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_9_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_213_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1);
  assign layer4_out_conc_213_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_213_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_10_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_215_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1);
  assign layer4_out_conc_215_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_215_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_11_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_217_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1);
  assign layer4_out_conc_217_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_217_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_12_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_219_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1);
  assign layer4_out_conc_219_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_219_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_13_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_221_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1);
  assign layer4_out_conc_221_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_221_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_14_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_223_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1);
  assign layer4_out_conc_223_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_223_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_15_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_225_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1);
  assign layer4_out_conc_225_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_225_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_16_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_227_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1);
  assign layer4_out_conc_227_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_227_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_17_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_229_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1);
  assign layer4_out_conc_229_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_229_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_18_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_231_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1);
  assign layer4_out_conc_231_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_231_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_19_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_233_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1);
  assign layer4_out_conc_233_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_233_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_20_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_235_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1);
  assign layer4_out_conc_235_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_235_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_21_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_237_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1);
  assign layer4_out_conc_237_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_237_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_22_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_239_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1);
  assign layer4_out_conc_239_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_239_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_23_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_241_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1);
  assign layer4_out_conc_241_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_241_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_24_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_243_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1);
  assign layer4_out_conc_243_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_243_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_25_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_245_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1);
  assign layer4_out_conc_245_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_245_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_26_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_247_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1);
  assign layer4_out_conc_247_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_247_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_27_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_249_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1);
  assign layer4_out_conc_249_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_249_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_28_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_251_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1);
  assign layer4_out_conc_251_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_251_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_29_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_253_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1);
  assign layer4_out_conc_253_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_253_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_30_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_255_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1);
  assign layer4_out_conc_255_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_255_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_31_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_257_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1);
  assign layer4_out_conc_257_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_257_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_32_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_259_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1);
  assign layer4_out_conc_259_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_259_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_33_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_261_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1);
  assign layer4_out_conc_261_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_261_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_34_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_263_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1);
  assign layer4_out_conc_263_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_263_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_35_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_265_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1);
  assign layer4_out_conc_265_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_265_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_36_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_267_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1);
  assign layer4_out_conc_267_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_267_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_37_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_269_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1);
  assign layer4_out_conc_269_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_269_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_38_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_271_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1);
  assign layer4_out_conc_271_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_271_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_39_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_273_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1);
  assign layer4_out_conc_273_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_273_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_40_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_275_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1);
  assign layer4_out_conc_275_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_275_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_41_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_277_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1);
  assign layer4_out_conc_277_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_277_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_42_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_279_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1);
  assign layer4_out_conc_279_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_279_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_43_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_281_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1);
  assign layer4_out_conc_281_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_281_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_44_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_283_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1);
  assign layer4_out_conc_283_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_283_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_45_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_285_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1);
  assign layer4_out_conc_285_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_285_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_46_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_287_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1);
  assign layer4_out_conc_287_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_287_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_47_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_289_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1);
  assign layer4_out_conc_289_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_289_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_48_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_291_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1);
  assign layer4_out_conc_291_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_291_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_49_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_293_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1);
  assign layer4_out_conc_293_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_293_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_50_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_295_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1);
  assign layer4_out_conc_295_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_295_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_51_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_297_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1);
  assign layer4_out_conc_297_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_297_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_52_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_299_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1);
  assign layer4_out_conc_299_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_299_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_53_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_301_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1);
  assign layer4_out_conc_301_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_301_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_54_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_303_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1);
  assign layer4_out_conc_303_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_303_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_55_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_305_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1);
  assign layer4_out_conc_305_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_305_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_56_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_307_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1);
  assign layer4_out_conc_307_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_307_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_57_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_309_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1);
  assign layer4_out_conc_309_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_309_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_58_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_311_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1);
  assign layer4_out_conc_311_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_311_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_59_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_313_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1);
  assign layer4_out_conc_313_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_313_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_60_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_315_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1);
  assign layer4_out_conc_315_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_315_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_61_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_317_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1);
  assign layer4_out_conc_317_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_317_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_62_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign layer4_out_conc_319_9 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[8:1]),
      8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1);
  assign layer4_out_conc_319_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign layer4_out_conc_319_0 = ((nnet_dense_latency_input_t_layer2_t_config2_acc_63_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9 = ((Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_0 = ((Accum1_14_Accum2_65_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9 = ((Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_0 = ((Accum1_14_Accum2_66_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9 = ((Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_0 = ((Accum1_14_Accum2_67_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9 = ((Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_0 = ((Accum1_14_Accum2_68_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9 = ((Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_0 = ((Accum1_14_Accum2_69_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9 = ((Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_0 = ((Accum1_14_Accum2_70_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9 = ((Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_0 = ((Accum1_14_Accum2_71_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9 = ((Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_0 = ((Accum1_14_Accum2_72_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9 = ((Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_0 = ((Accum1_14_Accum2_73_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9 = ((Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_0 = ((Accum1_14_Accum2_74_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9 = ((Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_0 = ((Accum1_14_Accum2_75_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9 = ((Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_0 = ((Accum1_14_Accum2_76_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9 = ((Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_0 = ((Accum1_14_Accum2_77_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_9 = ((Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_0 = ((Accum1_14_Accum2_78_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_9 = ((Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_0 = ((Accum1_14_Accum2_79_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_9 = ((Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_0 = ((Accum1_14_Accum2_80_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_9 = ((Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_0 = ((Accum1_14_Accum2_81_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_9 = ((Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_0 = ((Accum1_14_Accum2_82_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_9 = ((Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_0 = ((Accum1_14_Accum2_83_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_9 = ((Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_0 = ((Accum1_14_Accum2_84_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_9 = ((Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_0 = ((Accum1_14_Accum2_85_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_9 = ((Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_0 = ((Accum1_14_Accum2_86_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_9 = ((Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_0 = ((Accum1_14_Accum2_87_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_9 = ((Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_0 = ((Accum1_14_Accum2_88_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_9 = ((Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_0 = ((Accum1_14_Accum2_89_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_9 = ((Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_0 = ((Accum1_14_Accum2_90_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_9 = ((Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_0 = ((Accum1_14_Accum2_91_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_9 = ((Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_0 = ((Accum1_14_Accum2_92_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_9 = ((Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_0 = ((Accum1_14_Accum2_93_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_9 = ((Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_0 = ((Accum1_14_Accum2_94_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_9 = ((Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_0 = ((Accum1_14_Accum2_95_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_9 = ((Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_0 = ((Accum1_14_Accum2_96_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_9 = ((Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_0 = ((Accum1_14_Accum2_97_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_9 = ((Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_0 = ((Accum1_14_Accum2_98_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_9 = ((Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_0 = ((Accum1_14_Accum2_99_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_9 = ((Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_0 = ((Accum1_14_Accum2_100_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_9 = ((Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_0 = ((Accum1_14_Accum2_101_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_9 = ((Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_0 = ((Accum1_14_Accum2_102_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_9 = ((Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_0 = ((Accum1_14_Accum2_103_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_9 = ((Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_0 = ((Accum1_14_Accum2_104_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_9 = ((Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[9])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[8:1]), 8'b11111111,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_0 = ((Accum1_14_Accum2_107_Accum2_acc_1_ncse_sva_1[0])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  always @(posedge clk) begin
    if ( rst ) begin
      layer6_out_rsci_idat_15_0 <= 16'b0000000000000000;
      layer6_out_rsci_idat_31_16 <= 16'b0000000000000000;
      layer6_out_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else begin
      layer6_out_rsci_idat_15_0 <= nl_layer6_out_rsci_idat_15_0[15:0];
      layer6_out_rsci_idat_31_16 <= nl_layer6_out_rsci_idat_31_16[15:0];
      layer6_out_rsci_idat_47_32 <= nl_layer6_out_rsci_idat_47_32[15:0];
    end
  end
  assign nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_307_9 , layer4_out_conc_307_8_1 ,
      layer4_out_conc_307_0})) * $signed((w5_rsci_idat[859:855]));
  assign Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_309_9 , layer4_out_conc_309_8_1 ,
      layer4_out_conc_309_0})) * $signed((w5_rsci_idat[874:870]));
  assign Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_311_9 , layer4_out_conc_311_8_1 ,
      layer4_out_conc_311_0})) * $signed((w5_rsci_idat[889:885]));
  assign Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_313_9 , layer4_out_conc_313_8_1 ,
      layer4_out_conc_313_0})) * $signed((w5_rsci_idat[904:900]));
  assign Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_90_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_0}))
      * $signed((w5_rsci_idat[1339:1335]));
  assign Product1_1_90_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_90_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_91_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_0}))
      * $signed((w5_rsci_idat[1354:1350]));
  assign Product1_1_91_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_91_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_92_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_0}))
      * $signed((w5_rsci_idat[1369:1365]));
  assign Product1_1_92_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_92_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_93_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_0}))
      * $signed((w5_rsci_idat[1384:1380]));
  assign Product1_1_93_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_93_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_94_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_0}))
      * $signed((w5_rsci_idat[1399:1395]));
  assign Product1_1_94_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_94_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_95_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_0}))
      * $signed((w5_rsci_idat[1414:1410]));
  assign Product1_1_95_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_95_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_96_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_0}))
      * $signed((w5_rsci_idat[1429:1425]));
  assign Product1_1_96_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_96_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_97_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_0}))
      * $signed((w5_rsci_idat[1444:1440]));
  assign Product1_1_97_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_97_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_78_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_0}))
      * $signed((w5_rsci_idat[1159:1155]));
  assign Product1_1_78_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_78_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_79_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_0}))
      * $signed((w5_rsci_idat[1174:1170]));
  assign Product1_1_79_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_79_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_74_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_0}))
      * $signed((w5_rsci_idat[1099:1095]));
  assign Product1_1_74_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_74_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_75_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_0}))
      * $signed((w5_rsci_idat[1114:1110]));
  assign Product1_1_75_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_75_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_76_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_0}))
      * $signed((w5_rsci_idat[1129:1125]));
  assign Product1_1_76_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_76_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_77_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_0}))
      * $signed((w5_rsci_idat[1144:1140]));
  assign Product1_1_77_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_77_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_0}))
      * $signed((w5_rsci_idat[1189:1185]));
  assign Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_81_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_0}))
      * $signed((w5_rsci_idat[1204:1200]));
  assign Product1_1_81_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_81_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_86_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_0}))
      * $signed((w5_rsci_idat[1279:1275]));
  assign Product1_1_86_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_86_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_87_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_0}))
      * $signed((w5_rsci_idat[1294:1290]));
  assign Product1_1_87_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_87_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_82_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_0}))
      * $signed((w5_rsci_idat[1219:1215]));
  assign Product1_1_82_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_82_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_83_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_0}))
      * $signed((w5_rsci_idat[1234:1230]));
  assign Product1_1_83_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_83_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_84_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_0}))
      * $signed((w5_rsci_idat[1249:1245]));
  assign Product1_1_84_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_84_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_85_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_0}))
      * $signed((w5_rsci_idat[1264:1260]));
  assign Product1_1_85_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_85_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_88_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_0}))
      * $signed((w5_rsci_idat[1309:1305]));
  assign Product1_1_88_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_88_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_89_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_0}))
      * $signed((w5_rsci_idat[1324:1320]));
  assign Product1_1_89_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_89_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_275_9 , layer4_out_conc_275_8_1 ,
      layer4_out_conc_275_0})) * $signed((w5_rsci_idat[619:615]));
  assign Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_277_9 , layer4_out_conc_277_8_1 ,
      layer4_out_conc_277_0})) * $signed((w5_rsci_idat[634:630]));
  assign Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_279_9 , layer4_out_conc_279_8_1 ,
      layer4_out_conc_279_0})) * $signed((w5_rsci_idat[649:645]));
  assign Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_281_9 , layer4_out_conc_281_8_1 ,
      layer4_out_conc_281_0})) * $signed((w5_rsci_idat[664:660]));
  assign Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_283_9 , layer4_out_conc_283_8_1 ,
      layer4_out_conc_283_0})) * $signed((w5_rsci_idat[679:675]));
  assign Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_285_9 , layer4_out_conc_285_8_1 ,
      layer4_out_conc_285_0})) * $signed((w5_rsci_idat[694:690]));
  assign Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_287_9 , layer4_out_conc_287_8_1 ,
      layer4_out_conc_287_0})) * $signed((w5_rsci_idat[709:705]));
  assign Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_289_9 , layer4_out_conc_289_8_1 ,
      layer4_out_conc_289_0})) * $signed((w5_rsci_idat[724:720]));
  assign Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_299_9 , layer4_out_conc_299_8_1 ,
      layer4_out_conc_299_0})) * $signed((w5_rsci_idat[799:795]));
  assign Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_301_9 , layer4_out_conc_301_8_1 ,
      layer4_out_conc_301_0})) * $signed((w5_rsci_idat[814:810]));
  assign Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_303_9 , layer4_out_conc_303_8_1 ,
      layer4_out_conc_303_0})) * $signed((w5_rsci_idat[829:825]));
  assign Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_305_9 , layer4_out_conc_305_8_1 ,
      layer4_out_conc_305_0})) * $signed((w5_rsci_idat[844:840]));
  assign Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_291_9 , layer4_out_conc_291_8_1 ,
      layer4_out_conc_291_0})) * $signed((w5_rsci_idat[739:735]));
  assign Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_293_9 , layer4_out_conc_293_8_1 ,
      layer4_out_conc_293_0})) * $signed((w5_rsci_idat[754:750]));
  assign Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_295_9 , layer4_out_conc_295_8_1 ,
      layer4_out_conc_295_0})) * $signed((w5_rsci_idat[769:765]));
  assign Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_297_9 , layer4_out_conc_297_8_1 ,
      layer4_out_conc_297_0})) * $signed((w5_rsci_idat[784:780]));
  assign Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_315_9 , layer4_out_conc_315_8_1 ,
      layer4_out_conc_315_0})) * $signed((w5_rsci_idat[919:915]));
  assign Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_317_9 , layer4_out_conc_317_8_1 ,
      layer4_out_conc_317_0})) * $signed((w5_rsci_idat[934:930]));
  assign Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_319_9 , layer4_out_conc_319_8_1 ,
      layer4_out_conc_319_0})) * $signed((w5_rsci_idat[949:945]));
  assign Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_65_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_0}))
      * $signed((w5_rsci_idat[964:960]));
  assign Product1_1_65_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_65_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_70_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_0}))
      * $signed((w5_rsci_idat[1039:1035]));
  assign Product1_1_70_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_70_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_71_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_0}))
      * $signed((w5_rsci_idat[1054:1050]));
  assign Product1_1_71_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_71_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_72_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_0}))
      * $signed((w5_rsci_idat[1069:1065]));
  assign Product1_1_72_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_72_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_73_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_0}))
      * $signed((w5_rsci_idat[1084:1080]));
  assign Product1_1_73_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_73_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_66_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_0}))
      * $signed((w5_rsci_idat[979:975]));
  assign Product1_1_66_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_66_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_67_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_0}))
      * $signed((w5_rsci_idat[994:990]));
  assign Product1_1_67_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_67_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_68_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_0}))
      * $signed((w5_rsci_idat[1009:1005]));
  assign Product1_1_68_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_68_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_69_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_0}))
      * $signed((w5_rsci_idat[1024:1020]));
  assign Product1_1_69_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_69_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_102_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_0}))
      * $signed((w5_rsci_idat[1519:1515]));
  assign Product1_1_102_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_102_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_103_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_0}))
      * $signed((w5_rsci_idat[1534:1530]));
  assign Product1_1_103_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_103_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_104_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_0}))
      * $signed((w5_rsci_idat[1549:1545]));
  assign Product1_1_104_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_104_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_105_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_0}))
      * $signed((w5_rsci_idat[1564:1560]));
  assign Product1_1_105_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_105_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_98_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_0}))
      * $signed((w5_rsci_idat[1459:1455]));
  assign Product1_1_98_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_98_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_99_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_0}))
      * $signed((w5_rsci_idat[1474:1470]));
  assign Product1_1_99_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_99_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_100_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_0}))
      * $signed((w5_rsci_idat[1489:1485]));
  assign Product1_1_100_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_100_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_101_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_0}))
      * $signed((w5_rsci_idat[1504:1500]));
  assign Product1_1_101_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_101_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_386_nl = conv_s2s_11_16(readslicef_15_11_4(Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_90_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_91_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_92_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_93_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_94_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_95_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_96_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_97_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_78_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_79_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_74_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_75_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_76_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_77_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_80_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_81_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_86_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_87_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_82_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_83_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_84_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_85_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_88_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_89_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_65_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_70_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_71_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_72_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_73_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_66_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_67_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_68_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_69_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_102_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_103_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_104_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_105_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_98_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_99_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_100_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_101_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign Accum2_1_acc_386_nl = nl_Accum2_1_acc_386_nl[15:0];
  assign nl_Product1_1_126_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_0}))
      * $signed((w5_rsci_idat[1879:1875]));
  assign Product1_1_126_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_126_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_123_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_0}))
      * $signed((w5_rsci_idat[1834:1830]));
  assign Product1_1_123_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_123_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_118_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_0}))
      * $signed((w5_rsci_idat[1759:1755]));
  assign Product1_1_118_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_118_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_115_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_0}))
      * $signed((w5_rsci_idat[1714:1710]));
  assign Product1_1_115_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_115_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_122_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_0}))
      * $signed((w5_rsci_idat[1819:1815]));
  assign Product1_1_122_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_122_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_119_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_0}))
      * $signed((w5_rsci_idat[1774:1770]));
  assign Product1_1_119_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_119_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_203_9 , layer4_out_conc_203_8_1 ,
      layer4_out_conc_203_0})) * $signed((w5_rsci_idat[79:75]));
  assign Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_205_9 , layer4_out_conc_205_8_1 ,
      layer4_out_conc_205_0})) * $signed((w5_rsci_idat[94:90]));
  assign Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_195_9 , layer4_out_conc_195_8_1 ,
      layer4_out_conc_195_0})) * $signed((w5_rsci_idat[19:15]));
  assign Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_197_9 , layer4_out_conc_197_8_1 ,
      layer4_out_conc_197_0})) * $signed((w5_rsci_idat[34:30]));
  assign Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_199_9 , layer4_out_conc_199_8_1 ,
      layer4_out_conc_199_0})) * $signed((w5_rsci_idat[49:45]));
  assign Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_201_9 , layer4_out_conc_201_8_1 ,
      layer4_out_conc_201_0})) * $signed((w5_rsci_idat[64:60]));
  assign Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_114_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_0}))
      * $signed((w5_rsci_idat[1699:1695]));
  assign Product1_1_114_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_114_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_111_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_0}))
      * $signed((w5_rsci_idat[1654:1650]));
  assign Product1_1_111_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_111_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_112_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_0}))
      * $signed((w5_rsci_idat[1669:1665]));
  assign Product1_1_112_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_112_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_109_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_0}))
      * $signed((w5_rsci_idat[1624:1620]));
  assign Product1_1_109_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_109_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_389_nl = conv_s2s_5_6(b5_rsci_idat[4:0]) + conv_s2s_5_6(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1[10:6]);
  assign Accum2_1_acc_389_nl = nl_Accum2_1_acc_389_nl[5:0];
  assign nl_Product1_1_110_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_0}))
      * $signed((w5_rsci_idat[1639:1635]));
  assign Product1_1_110_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_110_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_108_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_0}))
      * $signed((w5_rsci_idat[1609:1605]));
  assign Product1_1_108_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_108_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_127_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_0}))
      * $signed((w5_rsci_idat[1894:1890]));
  assign Product1_1_127_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_127_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_106_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_0}))
      * $signed((w5_rsci_idat[1579:1575]));
  assign Product1_1_106_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_106_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_107_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_0}))
      * $signed((w5_rsci_idat[1594:1590]));
  assign Product1_1_107_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_107_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_128_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_0}))
      * $signed((w5_rsci_idat[1909:1905]));
  assign Product1_1_128_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_128_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_125_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_0}))
      * $signed((w5_rsci_idat[1864:1860]));
  assign Product1_1_125_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_125_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_124_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_0}))
      * $signed((w5_rsci_idat[1849:1845]));
  assign Product1_1_124_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_124_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_121_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_0}))
      * $signed((w5_rsci_idat[1804:1800]));
  assign Product1_1_121_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_121_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_120_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_0}))
      * $signed((w5_rsci_idat[1789:1785]));
  assign Product1_1_120_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_120_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_117_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_0}))
      * $signed((w5_rsci_idat[1744:1740]));
  assign Product1_1_117_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_117_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_116_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_0}))
      * $signed((w5_rsci_idat[1729:1725]));
  assign Product1_1_116_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_116_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_113_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_0}))
      * $signed((w5_rsci_idat[1684:1680]));
  assign Product1_1_113_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_113_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_207_9 , layer4_out_conc_207_8_1 ,
      layer4_out_conc_207_0})) * $signed((w5_rsci_idat[109:105]));
  assign Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_209_9 , layer4_out_conc_209_8_1 ,
      layer4_out_conc_209_0})) * $signed((w5_rsci_idat[124:120]));
  assign Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_385_nl = conv_s2s_11_16(readslicef_15_11_4(Product1_1_126_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_123_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_118_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_115_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_122_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_119_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_114_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_111_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_112_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_109_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_12_16({Accum2_1_acc_389_nl , (Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1[5:0])})
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_110_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_108_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_127_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_106_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_107_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_128_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_125_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_124_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_121_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_120_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_117_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_116_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_113_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign Accum2_1_acc_385_nl = nl_Accum2_1_acc_385_nl[15:0];
  assign nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_219_9 , layer4_out_conc_219_8_1 ,
      layer4_out_conc_219_0})) * $signed((w5_rsci_idat[199:195]));
  assign Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_221_9 , layer4_out_conc_221_8_1 ,
      layer4_out_conc_221_0})) * $signed((w5_rsci_idat[214:210]));
  assign Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_211_9 , layer4_out_conc_211_8_1 ,
      layer4_out_conc_211_0})) * $signed((w5_rsci_idat[139:135]));
  assign Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_213_9 , layer4_out_conc_213_8_1 ,
      layer4_out_conc_213_0})) * $signed((w5_rsci_idat[154:150]));
  assign Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_235_9 , layer4_out_conc_235_8_1 ,
      layer4_out_conc_235_0})) * $signed((w5_rsci_idat[319:315]));
  assign Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_237_9 , layer4_out_conc_237_8_1 ,
      layer4_out_conc_237_0})) * $signed((w5_rsci_idat[334:330]));
  assign Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_227_9 , layer4_out_conc_227_8_1 ,
      layer4_out_conc_227_0})) * $signed((w5_rsci_idat[259:255]));
  assign Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_229_9 , layer4_out_conc_229_8_1 ,
      layer4_out_conc_229_0})) * $signed((w5_rsci_idat[274:270]));
  assign Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_231_9 , layer4_out_conc_231_8_1 ,
      layer4_out_conc_231_0})) * $signed((w5_rsci_idat[289:285]));
  assign Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_233_9 , layer4_out_conc_233_8_1 ,
      layer4_out_conc_233_0})) * $signed((w5_rsci_idat[304:300]));
  assign Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_243_9 , layer4_out_conc_243_8_1 ,
      layer4_out_conc_243_0})) * $signed((w5_rsci_idat[379:375]));
  assign Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_245_9 , layer4_out_conc_245_8_1 ,
      layer4_out_conc_245_0})) * $signed((w5_rsci_idat[394:390]));
  assign Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_247_9 , layer4_out_conc_247_8_1 ,
      layer4_out_conc_247_0})) * $signed((w5_rsci_idat[409:405]));
  assign Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_249_9 , layer4_out_conc_249_8_1 ,
      layer4_out_conc_249_0})) * $signed((w5_rsci_idat[424:420]));
  assign Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_251_9 , layer4_out_conc_251_8_1 ,
      layer4_out_conc_251_0})) * $signed((w5_rsci_idat[439:435]));
  assign Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_253_9 , layer4_out_conc_253_8_1 ,
      layer4_out_conc_253_0})) * $signed((w5_rsci_idat[454:450]));
  assign Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_255_9 , layer4_out_conc_255_8_1 ,
      layer4_out_conc_255_0})) * $signed((w5_rsci_idat[469:465]));
  assign Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_257_9 , layer4_out_conc_257_8_1 ,
      layer4_out_conc_257_0})) * $signed((w5_rsci_idat[484:480]));
  assign Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_267_9 , layer4_out_conc_267_8_1 ,
      layer4_out_conc_267_0})) * $signed((w5_rsci_idat[559:555]));
  assign Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_269_9 , layer4_out_conc_269_8_1 ,
      layer4_out_conc_269_0})) * $signed((w5_rsci_idat[574:570]));
  assign Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_271_9 , layer4_out_conc_271_8_1 ,
      layer4_out_conc_271_0})) * $signed((w5_rsci_idat[589:585]));
  assign Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_273_9 , layer4_out_conc_273_8_1 ,
      layer4_out_conc_273_0})) * $signed((w5_rsci_idat[604:600]));
  assign Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_259_9 , layer4_out_conc_259_8_1 ,
      layer4_out_conc_259_0})) * $signed((w5_rsci_idat[499:495]));
  assign Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_261_9 , layer4_out_conc_261_8_1 ,
      layer4_out_conc_261_0})) * $signed((w5_rsci_idat[514:510]));
  assign Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_263_9 , layer4_out_conc_263_8_1 ,
      layer4_out_conc_263_0})) * $signed((w5_rsci_idat[529:525]));
  assign Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_265_9 , layer4_out_conc_265_8_1 ,
      layer4_out_conc_265_0})) * $signed((w5_rsci_idat[544:540]));
  assign Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_215_9 , layer4_out_conc_215_8_1 ,
      layer4_out_conc_215_0})) * $signed((w5_rsci_idat[169:165]));
  assign Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_217_9 , layer4_out_conc_217_8_1 ,
      layer4_out_conc_217_0})) * $signed((w5_rsci_idat[184:180]));
  assign Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_223_9 , layer4_out_conc_223_8_1 ,
      layer4_out_conc_223_0})) * $signed((w5_rsci_idat[229:225]));
  assign Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_225_9 , layer4_out_conc_225_8_1 ,
      layer4_out_conc_225_0})) * $signed((w5_rsci_idat[244:240]));
  assign Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_239_9 , layer4_out_conc_239_8_1 ,
      layer4_out_conc_239_0})) * $signed((w5_rsci_idat[349:345]));
  assign Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_241_9 , layer4_out_conc_241_8_1 ,
      layer4_out_conc_241_0})) * $signed((w5_rsci_idat[364:360]));
  assign Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_layer6_out_rsci_idat_15_0  = Accum2_1_acc_386_nl + Accum2_1_acc_385_nl
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_307_9 , layer4_out_conc_307_8_1 ,
      layer4_out_conc_307_0})) * $signed((w5_rsci_idat[864:860]));
  assign Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_309_9 , layer4_out_conc_309_8_1 ,
      layer4_out_conc_309_0})) * $signed((w5_rsci_idat[879:875]));
  assign Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_311_9 , layer4_out_conc_311_8_1 ,
      layer4_out_conc_311_0})) * $signed((w5_rsci_idat[894:890]));
  assign Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_313_9 , layer4_out_conc_313_8_1 ,
      layer4_out_conc_313_0})) * $signed((w5_rsci_idat[909:905]));
  assign Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_90_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_0}))
      * $signed((w5_rsci_idat[1344:1340]));
  assign Product1_1_90_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_90_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_91_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_0}))
      * $signed((w5_rsci_idat[1359:1355]));
  assign Product1_1_91_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_91_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_92_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_0}))
      * $signed((w5_rsci_idat[1374:1370]));
  assign Product1_1_92_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_92_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_93_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_0}))
      * $signed((w5_rsci_idat[1389:1385]));
  assign Product1_1_93_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_93_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_94_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_0}))
      * $signed((w5_rsci_idat[1404:1400]));
  assign Product1_1_94_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_94_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_95_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_0}))
      * $signed((w5_rsci_idat[1419:1415]));
  assign Product1_1_95_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_95_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_96_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_0}))
      * $signed((w5_rsci_idat[1434:1430]));
  assign Product1_1_96_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_96_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_97_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_0}))
      * $signed((w5_rsci_idat[1449:1445]));
  assign Product1_1_97_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_97_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_78_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_0}))
      * $signed((w5_rsci_idat[1164:1160]));
  assign Product1_1_78_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_78_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_79_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_0}))
      * $signed((w5_rsci_idat[1179:1175]));
  assign Product1_1_79_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_79_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_74_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_0}))
      * $signed((w5_rsci_idat[1104:1100]));
  assign Product1_1_74_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_74_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_75_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_0}))
      * $signed((w5_rsci_idat[1119:1115]));
  assign Product1_1_75_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_75_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_76_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_0}))
      * $signed((w5_rsci_idat[1134:1130]));
  assign Product1_1_76_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_76_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_77_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_0}))
      * $signed((w5_rsci_idat[1149:1145]));
  assign Product1_1_77_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_77_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_80_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_0}))
      * $signed((w5_rsci_idat[1194:1190]));
  assign Product1_1_80_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_80_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_81_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_0}))
      * $signed((w5_rsci_idat[1209:1205]));
  assign Product1_1_81_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_81_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_86_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_0}))
      * $signed((w5_rsci_idat[1284:1280]));
  assign Product1_1_86_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_86_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_87_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_0}))
      * $signed((w5_rsci_idat[1299:1295]));
  assign Product1_1_87_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_87_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_82_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_0}))
      * $signed((w5_rsci_idat[1224:1220]));
  assign Product1_1_82_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_82_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_83_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_0}))
      * $signed((w5_rsci_idat[1239:1235]));
  assign Product1_1_83_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_83_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_84_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_0}))
      * $signed((w5_rsci_idat[1254:1250]));
  assign Product1_1_84_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_84_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_85_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_0}))
      * $signed((w5_rsci_idat[1269:1265]));
  assign Product1_1_85_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_85_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_88_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_0}))
      * $signed((w5_rsci_idat[1314:1310]));
  assign Product1_1_88_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_88_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_89_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_0}))
      * $signed((w5_rsci_idat[1329:1325]));
  assign Product1_1_89_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_89_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_275_9 , layer4_out_conc_275_8_1 ,
      layer4_out_conc_275_0})) * $signed((w5_rsci_idat[624:620]));
  assign Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_277_9 , layer4_out_conc_277_8_1 ,
      layer4_out_conc_277_0})) * $signed((w5_rsci_idat[639:635]));
  assign Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_279_9 , layer4_out_conc_279_8_1 ,
      layer4_out_conc_279_0})) * $signed((w5_rsci_idat[654:650]));
  assign Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_281_9 , layer4_out_conc_281_8_1 ,
      layer4_out_conc_281_0})) * $signed((w5_rsci_idat[669:665]));
  assign Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_283_9 , layer4_out_conc_283_8_1 ,
      layer4_out_conc_283_0})) * $signed((w5_rsci_idat[684:680]));
  assign Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_285_9 , layer4_out_conc_285_8_1 ,
      layer4_out_conc_285_0})) * $signed((w5_rsci_idat[699:695]));
  assign Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_287_9 , layer4_out_conc_287_8_1 ,
      layer4_out_conc_287_0})) * $signed((w5_rsci_idat[714:710]));
  assign Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_289_9 , layer4_out_conc_289_8_1 ,
      layer4_out_conc_289_0})) * $signed((w5_rsci_idat[729:725]));
  assign Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_299_9 , layer4_out_conc_299_8_1 ,
      layer4_out_conc_299_0})) * $signed((w5_rsci_idat[804:800]));
  assign Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_301_9 , layer4_out_conc_301_8_1 ,
      layer4_out_conc_301_0})) * $signed((w5_rsci_idat[819:815]));
  assign Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_303_9 , layer4_out_conc_303_8_1 ,
      layer4_out_conc_303_0})) * $signed((w5_rsci_idat[834:830]));
  assign Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_305_9 , layer4_out_conc_305_8_1 ,
      layer4_out_conc_305_0})) * $signed((w5_rsci_idat[849:845]));
  assign Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_291_9 , layer4_out_conc_291_8_1 ,
      layer4_out_conc_291_0})) * $signed((w5_rsci_idat[744:740]));
  assign Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_293_9 , layer4_out_conc_293_8_1 ,
      layer4_out_conc_293_0})) * $signed((w5_rsci_idat[759:755]));
  assign Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_295_9 , layer4_out_conc_295_8_1 ,
      layer4_out_conc_295_0})) * $signed((w5_rsci_idat[774:770]));
  assign Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_297_9 , layer4_out_conc_297_8_1 ,
      layer4_out_conc_297_0})) * $signed((w5_rsci_idat[789:785]));
  assign Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_315_9 , layer4_out_conc_315_8_1 ,
      layer4_out_conc_315_0})) * $signed((w5_rsci_idat[924:920]));
  assign Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_317_9 , layer4_out_conc_317_8_1 ,
      layer4_out_conc_317_0})) * $signed((w5_rsci_idat[939:935]));
  assign Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_319_9 , layer4_out_conc_319_8_1 ,
      layer4_out_conc_319_0})) * $signed((w5_rsci_idat[954:950]));
  assign Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_65_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_0}))
      * $signed((w5_rsci_idat[969:965]));
  assign Product1_1_65_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_65_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_70_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_0}))
      * $signed((w5_rsci_idat[1044:1040]));
  assign Product1_1_70_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_70_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_71_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_0}))
      * $signed((w5_rsci_idat[1059:1055]));
  assign Product1_1_71_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_71_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_72_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_0}))
      * $signed((w5_rsci_idat[1074:1070]));
  assign Product1_1_72_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_72_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_73_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_0}))
      * $signed((w5_rsci_idat[1089:1085]));
  assign Product1_1_73_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_73_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_66_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_0}))
      * $signed((w5_rsci_idat[984:980]));
  assign Product1_1_66_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_66_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_67_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_0}))
      * $signed((w5_rsci_idat[999:995]));
  assign Product1_1_67_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_67_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_68_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_0}))
      * $signed((w5_rsci_idat[1014:1010]));
  assign Product1_1_68_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_68_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_69_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_0}))
      * $signed((w5_rsci_idat[1029:1025]));
  assign Product1_1_69_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_69_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_102_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_0}))
      * $signed((w5_rsci_idat[1524:1520]));
  assign Product1_1_102_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_102_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_103_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_0}))
      * $signed((w5_rsci_idat[1539:1535]));
  assign Product1_1_103_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_103_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_104_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_0}))
      * $signed((w5_rsci_idat[1554:1550]));
  assign Product1_1_104_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_104_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_105_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_0}))
      * $signed((w5_rsci_idat[1569:1565]));
  assign Product1_1_105_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_105_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_98_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_0}))
      * $signed((w5_rsci_idat[1464:1460]));
  assign Product1_1_98_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_98_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_99_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_0}))
      * $signed((w5_rsci_idat[1479:1475]));
  assign Product1_1_99_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_99_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_100_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_0}))
      * $signed((w5_rsci_idat[1494:1490]));
  assign Product1_1_100_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_100_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_101_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_0}))
      * $signed((w5_rsci_idat[1509:1505]));
  assign Product1_1_101_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_101_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_259_nl = conv_s2s_11_16(readslicef_15_11_4(Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_90_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_91_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_92_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_93_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_94_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_95_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_96_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_97_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_78_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_79_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_74_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_75_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_76_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_77_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_80_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_81_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_86_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_87_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_82_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_83_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_84_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_85_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_88_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_89_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_65_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_70_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_71_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_72_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_73_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_66_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_67_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_68_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_69_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_102_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_103_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_104_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_105_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_98_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_99_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_100_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_101_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign Accum2_1_acc_259_nl = nl_Accum2_1_acc_259_nl[15:0];
  assign nl_Product1_1_126_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_0}))
      * $signed((w5_rsci_idat[1884:1880]));
  assign Product1_1_126_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_126_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_123_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_0}))
      * $signed((w5_rsci_idat[1839:1835]));
  assign Product1_1_123_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_123_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_118_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_0}))
      * $signed((w5_rsci_idat[1764:1760]));
  assign Product1_1_118_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_118_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_115_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_0}))
      * $signed((w5_rsci_idat[1719:1715]));
  assign Product1_1_115_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_115_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_122_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_0}))
      * $signed((w5_rsci_idat[1824:1820]));
  assign Product1_1_122_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_122_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_119_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_0}))
      * $signed((w5_rsci_idat[1779:1775]));
  assign Product1_1_119_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_119_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_203_9 , layer4_out_conc_203_8_1 ,
      layer4_out_conc_203_0})) * $signed((w5_rsci_idat[84:80]));
  assign Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_205_9 , layer4_out_conc_205_8_1 ,
      layer4_out_conc_205_0})) * $signed((w5_rsci_idat[99:95]));
  assign Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_195_9 , layer4_out_conc_195_8_1 ,
      layer4_out_conc_195_0})) * $signed((w5_rsci_idat[24:20]));
  assign Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_197_9 , layer4_out_conc_197_8_1 ,
      layer4_out_conc_197_0})) * $signed((w5_rsci_idat[39:35]));
  assign Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_199_9 , layer4_out_conc_199_8_1 ,
      layer4_out_conc_199_0})) * $signed((w5_rsci_idat[54:50]));
  assign Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_201_9 , layer4_out_conc_201_8_1 ,
      layer4_out_conc_201_0})) * $signed((w5_rsci_idat[69:65]));
  assign Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_114_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_0}))
      * $signed((w5_rsci_idat[1704:1700]));
  assign Product1_1_114_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_114_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_111_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_0}))
      * $signed((w5_rsci_idat[1659:1655]));
  assign Product1_1_111_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_111_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_112_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_0}))
      * $signed((w5_rsci_idat[1674:1670]));
  assign Product1_1_112_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_112_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_109_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_0}))
      * $signed((w5_rsci_idat[1629:1625]));
  assign Product1_1_109_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_109_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_388_nl = conv_s2s_5_6(b5_rsci_idat[9:5]) + conv_s2s_5_6(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1[10:6]);
  assign Accum2_1_acc_388_nl = nl_Accum2_1_acc_388_nl[5:0];
  assign nl_Product1_1_110_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_0}))
      * $signed((w5_rsci_idat[1644:1640]));
  assign Product1_1_110_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_110_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_108_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_0}))
      * $signed((w5_rsci_idat[1614:1610]));
  assign Product1_1_108_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_108_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_127_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_0}))
      * $signed((w5_rsci_idat[1899:1895]));
  assign Product1_1_127_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_127_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_106_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_0}))
      * $signed((w5_rsci_idat[1584:1580]));
  assign Product1_1_106_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_106_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_107_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_384_0}))
      * $signed((w5_rsci_idat[1599:1595]));
  assign Product1_1_107_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_107_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_128_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_0}))
      * $signed((w5_rsci_idat[1914:1910]));
  assign Product1_1_128_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_128_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_125_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_0}))
      * $signed((w5_rsci_idat[1869:1865]));
  assign Product1_1_125_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_125_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_124_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_0}))
      * $signed((w5_rsci_idat[1854:1850]));
  assign Product1_1_124_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_124_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_121_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_0}))
      * $signed((w5_rsci_idat[1809:1805]));
  assign Product1_1_121_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_121_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_120_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_0}))
      * $signed((w5_rsci_idat[1794:1790]));
  assign Product1_1_120_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_120_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_117_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_0}))
      * $signed((w5_rsci_idat[1749:1745]));
  assign Product1_1_117_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_117_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_116_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_0}))
      * $signed((w5_rsci_idat[1734:1730]));
  assign Product1_1_116_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_116_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_113_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_0}))
      * $signed((w5_rsci_idat[1689:1685]));
  assign Product1_1_113_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_113_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_207_9 , layer4_out_conc_207_8_1 ,
      layer4_out_conc_207_0})) * $signed((w5_rsci_idat[114:110]));
  assign Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_209_9 , layer4_out_conc_209_8_1 ,
      layer4_out_conc_209_0})) * $signed((w5_rsci_idat[129:125]));
  assign Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_258_nl = conv_s2s_11_16(readslicef_15_11_4(Product1_1_126_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_123_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_118_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_115_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_122_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_119_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_114_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_111_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_112_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_109_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_12_16({Accum2_1_acc_388_nl , (Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1[5:0])})
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_110_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_108_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_127_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_106_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_107_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_128_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_125_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_124_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_121_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_120_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_117_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_116_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_113_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign Accum2_1_acc_258_nl = nl_Accum2_1_acc_258_nl[15:0];
  assign nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_219_9 , layer4_out_conc_219_8_1 ,
      layer4_out_conc_219_0})) * $signed((w5_rsci_idat[204:200]));
  assign Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_221_9 , layer4_out_conc_221_8_1 ,
      layer4_out_conc_221_0})) * $signed((w5_rsci_idat[219:215]));
  assign Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_211_9 , layer4_out_conc_211_8_1 ,
      layer4_out_conc_211_0})) * $signed((w5_rsci_idat[144:140]));
  assign Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_213_9 , layer4_out_conc_213_8_1 ,
      layer4_out_conc_213_0})) * $signed((w5_rsci_idat[159:155]));
  assign Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_235_9 , layer4_out_conc_235_8_1 ,
      layer4_out_conc_235_0})) * $signed((w5_rsci_idat[324:320]));
  assign Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_237_9 , layer4_out_conc_237_8_1 ,
      layer4_out_conc_237_0})) * $signed((w5_rsci_idat[339:335]));
  assign Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_227_9 , layer4_out_conc_227_8_1 ,
      layer4_out_conc_227_0})) * $signed((w5_rsci_idat[264:260]));
  assign Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_229_9 , layer4_out_conc_229_8_1 ,
      layer4_out_conc_229_0})) * $signed((w5_rsci_idat[279:275]));
  assign Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_231_9 , layer4_out_conc_231_8_1 ,
      layer4_out_conc_231_0})) * $signed((w5_rsci_idat[294:290]));
  assign Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_233_9 , layer4_out_conc_233_8_1 ,
      layer4_out_conc_233_0})) * $signed((w5_rsci_idat[309:305]));
  assign Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_243_9 , layer4_out_conc_243_8_1 ,
      layer4_out_conc_243_0})) * $signed((w5_rsci_idat[384:380]));
  assign Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_245_9 , layer4_out_conc_245_8_1 ,
      layer4_out_conc_245_0})) * $signed((w5_rsci_idat[399:395]));
  assign Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_247_9 , layer4_out_conc_247_8_1 ,
      layer4_out_conc_247_0})) * $signed((w5_rsci_idat[414:410]));
  assign Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_249_9 , layer4_out_conc_249_8_1 ,
      layer4_out_conc_249_0})) * $signed((w5_rsci_idat[429:425]));
  assign Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_251_9 , layer4_out_conc_251_8_1 ,
      layer4_out_conc_251_0})) * $signed((w5_rsci_idat[444:440]));
  assign Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_253_9 , layer4_out_conc_253_8_1 ,
      layer4_out_conc_253_0})) * $signed((w5_rsci_idat[459:455]));
  assign Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_255_9 , layer4_out_conc_255_8_1 ,
      layer4_out_conc_255_0})) * $signed((w5_rsci_idat[474:470]));
  assign Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_257_9 , layer4_out_conc_257_8_1 ,
      layer4_out_conc_257_0})) * $signed((w5_rsci_idat[489:485]));
  assign Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_267_9 , layer4_out_conc_267_8_1 ,
      layer4_out_conc_267_0})) * $signed((w5_rsci_idat[564:560]));
  assign Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_269_9 , layer4_out_conc_269_8_1 ,
      layer4_out_conc_269_0})) * $signed((w5_rsci_idat[579:575]));
  assign Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_271_9 , layer4_out_conc_271_8_1 ,
      layer4_out_conc_271_0})) * $signed((w5_rsci_idat[594:590]));
  assign Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_273_9 , layer4_out_conc_273_8_1 ,
      layer4_out_conc_273_0})) * $signed((w5_rsci_idat[609:605]));
  assign Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_259_9 , layer4_out_conc_259_8_1 ,
      layer4_out_conc_259_0})) * $signed((w5_rsci_idat[504:500]));
  assign Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_261_9 , layer4_out_conc_261_8_1 ,
      layer4_out_conc_261_0})) * $signed((w5_rsci_idat[519:515]));
  assign Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_263_9 , layer4_out_conc_263_8_1 ,
      layer4_out_conc_263_0})) * $signed((w5_rsci_idat[534:530]));
  assign Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_265_9 , layer4_out_conc_265_8_1 ,
      layer4_out_conc_265_0})) * $signed((w5_rsci_idat[549:545]));
  assign Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_215_9 , layer4_out_conc_215_8_1 ,
      layer4_out_conc_215_0})) * $signed((w5_rsci_idat[174:170]));
  assign Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_217_9 , layer4_out_conc_217_8_1 ,
      layer4_out_conc_217_0})) * $signed((w5_rsci_idat[189:185]));
  assign Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_223_9 , layer4_out_conc_223_8_1 ,
      layer4_out_conc_223_0})) * $signed((w5_rsci_idat[234:230]));
  assign Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_225_9 , layer4_out_conc_225_8_1 ,
      layer4_out_conc_225_0})) * $signed((w5_rsci_idat[249:245]));
  assign Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_239_9 , layer4_out_conc_239_8_1 ,
      layer4_out_conc_239_0})) * $signed((w5_rsci_idat[354:350]));
  assign Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_241_9 , layer4_out_conc_241_8_1 ,
      layer4_out_conc_241_0})) * $signed((w5_rsci_idat[369:365]));
  assign Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_layer6_out_rsci_idat_31_16  = Accum2_1_acc_259_nl + Accum2_1_acc_258_nl
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_305_9 , layer4_out_conc_305_8_1 ,
      layer4_out_conc_305_0})) * $signed((w5_rsci_idat[854:850]));
  assign Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_307_9 , layer4_out_conc_307_8_1 ,
      layer4_out_conc_307_0})) * $signed((w5_rsci_idat[869:865]));
  assign Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_309_9 , layer4_out_conc_309_8_1 ,
      layer4_out_conc_309_0})) * $signed((w5_rsci_idat[884:880]));
  assign Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_311_9 , layer4_out_conc_311_8_1 ,
      layer4_out_conc_311_0})) * $signed((w5_rsci_idat[899:895]));
  assign Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_89_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_352_0}))
      * $signed((w5_rsci_idat[1334:1330]));
  assign Product1_1_89_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_89_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_90_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_354_0}))
      * $signed((w5_rsci_idat[1349:1345]));
  assign Product1_1_90_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_90_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_91_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_356_0}))
      * $signed((w5_rsci_idat[1364:1360]));
  assign Product1_1_91_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_91_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_92_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_358_0}))
      * $signed((w5_rsci_idat[1379:1375]));
  assign Product1_1_92_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_92_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_93_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_360_0}))
      * $signed((w5_rsci_idat[1394:1390]));
  assign Product1_1_93_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_93_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_94_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_362_0}))
      * $signed((w5_rsci_idat[1409:1405]));
  assign Product1_1_94_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_94_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_95_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_364_0}))
      * $signed((w5_rsci_idat[1424:1420]));
  assign Product1_1_95_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_95_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_96_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_366_0}))
      * $signed((w5_rsci_idat[1439:1435]));
  assign Product1_1_96_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_96_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_77_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_0}))
      * $signed((w5_rsci_idat[1154:1150]));
  assign Product1_1_77_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_77_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_78_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_330_0}))
      * $signed((w5_rsci_idat[1169:1165]));
  assign Product1_1_78_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_78_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_73_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_0}))
      * $signed((w5_rsci_idat[1094:1090]));
  assign Product1_1_73_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_73_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_74_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_0}))
      * $signed((w5_rsci_idat[1109:1105]));
  assign Product1_1_74_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_74_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_75_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_0}))
      * $signed((w5_rsci_idat[1124:1120]));
  assign Product1_1_75_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_75_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_76_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_0}))
      * $signed((w5_rsci_idat[1139:1135]));
  assign Product1_1_76_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_76_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_79_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_332_0}))
      * $signed((w5_rsci_idat[1184:1180]));
  assign Product1_1_79_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_79_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_80_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_334_0}))
      * $signed((w5_rsci_idat[1199:1195]));
  assign Product1_1_80_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_80_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_85_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_344_0}))
      * $signed((w5_rsci_idat[1274:1270]));
  assign Product1_1_85_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_85_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_86_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_346_0}))
      * $signed((w5_rsci_idat[1289:1285]));
  assign Product1_1_86_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_86_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_81_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_336_0}))
      * $signed((w5_rsci_idat[1214:1210]));
  assign Product1_1_81_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_81_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_82_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_338_0}))
      * $signed((w5_rsci_idat[1229:1225]));
  assign Product1_1_82_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_82_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_83_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_340_0}))
      * $signed((w5_rsci_idat[1244:1240]));
  assign Product1_1_83_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_83_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_84_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_342_0}))
      * $signed((w5_rsci_idat[1259:1255]));
  assign Product1_1_84_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_84_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_87_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_348_0}))
      * $signed((w5_rsci_idat[1304:1300]));
  assign Product1_1_87_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_87_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_88_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_350_0}))
      * $signed((w5_rsci_idat[1319:1315]));
  assign Product1_1_88_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_88_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_273_9 , layer4_out_conc_273_8_1 ,
      layer4_out_conc_273_0})) * $signed((w5_rsci_idat[614:610]));
  assign Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_275_9 , layer4_out_conc_275_8_1 ,
      layer4_out_conc_275_0})) * $signed((w5_rsci_idat[629:625]));
  assign Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_277_9 , layer4_out_conc_277_8_1 ,
      layer4_out_conc_277_0})) * $signed((w5_rsci_idat[644:640]));
  assign Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_279_9 , layer4_out_conc_279_8_1 ,
      layer4_out_conc_279_0})) * $signed((w5_rsci_idat[659:655]));
  assign Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_281_9 , layer4_out_conc_281_8_1 ,
      layer4_out_conc_281_0})) * $signed((w5_rsci_idat[674:670]));
  assign Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_283_9 , layer4_out_conc_283_8_1 ,
      layer4_out_conc_283_0})) * $signed((w5_rsci_idat[689:685]));
  assign Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_285_9 , layer4_out_conc_285_8_1 ,
      layer4_out_conc_285_0})) * $signed((w5_rsci_idat[704:700]));
  assign Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_287_9 , layer4_out_conc_287_8_1 ,
      layer4_out_conc_287_0})) * $signed((w5_rsci_idat[719:715]));
  assign Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_297_9 , layer4_out_conc_297_8_1 ,
      layer4_out_conc_297_0})) * $signed((w5_rsci_idat[794:790]));
  assign Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_299_9 , layer4_out_conc_299_8_1 ,
      layer4_out_conc_299_0})) * $signed((w5_rsci_idat[809:805]));
  assign Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_301_9 , layer4_out_conc_301_8_1 ,
      layer4_out_conc_301_0})) * $signed((w5_rsci_idat[824:820]));
  assign Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_303_9 , layer4_out_conc_303_8_1 ,
      layer4_out_conc_303_0})) * $signed((w5_rsci_idat[839:835]));
  assign Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_289_9 , layer4_out_conc_289_8_1 ,
      layer4_out_conc_289_0})) * $signed((w5_rsci_idat[734:730]));
  assign Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_291_9 , layer4_out_conc_291_8_1 ,
      layer4_out_conc_291_0})) * $signed((w5_rsci_idat[749:745]));
  assign Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_293_9 , layer4_out_conc_293_8_1 ,
      layer4_out_conc_293_0})) * $signed((w5_rsci_idat[764:760]));
  assign Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_295_9 , layer4_out_conc_295_8_1 ,
      layer4_out_conc_295_0})) * $signed((w5_rsci_idat[779:775]));
  assign Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_313_9 , layer4_out_conc_313_8_1 ,
      layer4_out_conc_313_0})) * $signed((w5_rsci_idat[914:910]));
  assign Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_315_9 , layer4_out_conc_315_8_1 ,
      layer4_out_conc_315_0})) * $signed((w5_rsci_idat[929:925]));
  assign Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_317_9 , layer4_out_conc_317_8_1 ,
      layer4_out_conc_317_0})) * $signed((w5_rsci_idat[944:940]));
  assign Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_319_9 , layer4_out_conc_319_8_1 ,
      layer4_out_conc_319_0})) * $signed((w5_rsci_idat[959:955]));
  assign Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_69_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_0}))
      * $signed((w5_rsci_idat[1034:1030]));
  assign Product1_1_69_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_69_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_70_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_0}))
      * $signed((w5_rsci_idat[1049:1045]));
  assign Product1_1_70_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_70_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_71_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_0}))
      * $signed((w5_rsci_idat[1064:1060]));
  assign Product1_1_71_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_71_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_72_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_0}))
      * $signed((w5_rsci_idat[1079:1075]));
  assign Product1_1_72_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_72_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_65_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_0}))
      * $signed((w5_rsci_idat[974:970]));
  assign Product1_1_65_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_65_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_66_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_0}))
      * $signed((w5_rsci_idat[989:985]));
  assign Product1_1_66_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_66_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_67_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_0}))
      * $signed((w5_rsci_idat[1004:1000]));
  assign Product1_1_67_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_67_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_68_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_0}))
      * $signed((w5_rsci_idat[1019:1015]));
  assign Product1_1_68_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_68_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_101_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_376_0}))
      * $signed((w5_rsci_idat[1514:1510]));
  assign Product1_1_101_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_101_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_102_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_378_0}))
      * $signed((w5_rsci_idat[1529:1525]));
  assign Product1_1_102_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_102_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_103_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_380_0}))
      * $signed((w5_rsci_idat[1544:1540]));
  assign Product1_1_103_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_103_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_104_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_382_0}))
      * $signed((w5_rsci_idat[1559:1555]));
  assign Product1_1_104_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_104_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_97_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_368_0}))
      * $signed((w5_rsci_idat[1454:1450]));
  assign Product1_1_97_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_97_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_98_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_370_0}))
      * $signed((w5_rsci_idat[1469:1465]));
  assign Product1_1_98_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_98_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_99_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_372_0}))
      * $signed((w5_rsci_idat[1484:1480]));
  assign Product1_1_99_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_99_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_100_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_374_0}))
      * $signed((w5_rsci_idat[1499:1495]));
  assign Product1_1_100_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_100_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_132_nl = conv_s2s_11_16(readslicef_15_11_4(Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_89_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_90_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_91_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_92_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_93_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_94_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_95_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_96_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_77_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_78_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_73_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_74_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_75_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_76_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_79_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_80_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_85_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_86_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_81_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_82_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_83_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_84_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_87_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_88_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_69_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_70_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_71_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_72_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_65_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_66_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_67_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_68_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_101_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_102_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_103_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_104_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_97_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_98_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_99_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_100_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign Accum2_1_acc_132_nl = nl_Accum2_1_acc_132_nl[15:0];
  assign nl_Product1_1_124_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_0}))
      * $signed((w5_rsci_idat[1859:1855]));
  assign Product1_1_124_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_124_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_125_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_0}))
      * $signed((w5_rsci_idat[1874:1870]));
  assign Product1_1_125_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_125_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_116_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_0}))
      * $signed((w5_rsci_idat[1739:1735]));
  assign Product1_1_116_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_116_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_117_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_0}))
      * $signed((w5_rsci_idat[1754:1750]));
  assign Product1_1_117_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_117_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_120_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_0}))
      * $signed((w5_rsci_idat[1799:1795]));
  assign Product1_1_120_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_120_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_121_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_0}))
      * $signed((w5_rsci_idat[1814:1810]));
  assign Product1_1_121_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_121_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_201_9 , layer4_out_conc_201_8_1 ,
      layer4_out_conc_201_0})) * $signed((w5_rsci_idat[74:70]));
  assign Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_203_9 , layer4_out_conc_203_8_1 ,
      layer4_out_conc_203_0})) * $signed((w5_rsci_idat[89:85]));
  assign Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_193_9 , layer4_out_conc_193_8_1 ,
      layer4_out_conc_193_0})) * $signed((w5_rsci_idat[14:10]));
  assign Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_195_9 , layer4_out_conc_195_8_1 ,
      layer4_out_conc_195_0})) * $signed((w5_rsci_idat[29:25]));
  assign Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_197_9 , layer4_out_conc_197_8_1 ,
      layer4_out_conc_197_0})) * $signed((w5_rsci_idat[44:40]));
  assign Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_199_9 , layer4_out_conc_199_8_1 ,
      layer4_out_conc_199_0})) * $signed((w5_rsci_idat[59:55]));
  assign Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_112_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_0}))
      * $signed((w5_rsci_idat[1679:1675]));
  assign Product1_1_112_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_112_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_113_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_0}))
      * $signed((w5_rsci_idat[1694:1690]));
  assign Product1_1_113_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_113_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_110_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_0}))
      * $signed((w5_rsci_idat[1649:1645]));
  assign Product1_1_110_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_110_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_111_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_0}))
      * $signed((w5_rsci_idat[1664:1660]));
  assign Product1_1_111_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_111_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_390_nl = conv_s2s_5_6(Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1[10:6])
      + conv_s2s_5_6(b5_rsci_idat[14:10]);
  assign Accum2_1_acc_390_nl = nl_Accum2_1_acc_390_nl[5:0];
  assign nl_Product1_1_108_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_0}))
      * $signed((w5_rsci_idat[1619:1615]));
  assign Product1_1_108_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_108_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_109_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_0}))
      * $signed((w5_rsci_idat[1634:1630]));
  assign Product1_1_109_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_109_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_126_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_0}))
      * $signed((w5_rsci_idat[1889:1885]));
  assign Product1_1_126_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_126_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_105_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_0}))
      * $signed((w5_rsci_idat[1574:1570]));
  assign Product1_1_105_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_105_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_106_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_0}))
      * $signed((w5_rsci_idat[1589:1585]));
  assign Product1_1_106_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_106_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_127_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_0}))
      * $signed((w5_rsci_idat[1904:1900]));
  assign Product1_1_127_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_127_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_128_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_0}))
      * $signed((w5_rsci_idat[1919:1915]));
  assign Product1_1_128_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_128_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_122_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_0}))
      * $signed((w5_rsci_idat[1829:1825]));
  assign Product1_1_122_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_122_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_123_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_0}))
      * $signed((w5_rsci_idat[1844:1840]));
  assign Product1_1_123_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_123_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_118_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_0}))
      * $signed((w5_rsci_idat[1769:1765]));
  assign Product1_1_118_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_118_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_119_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_0}))
      * $signed((w5_rsci_idat[1784:1780]));
  assign Product1_1_119_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_119_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_114_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_0}))
      * $signed((w5_rsci_idat[1709:1705]));
  assign Product1_1_114_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_114_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_115_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_1 , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_0}))
      * $signed((w5_rsci_idat[1724:1720]));
  assign Product1_1_115_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_115_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_205_9 , layer4_out_conc_205_8_1 ,
      layer4_out_conc_205_0})) * $signed((w5_rsci_idat[104:100]));
  assign Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_207_9 , layer4_out_conc_207_8_1 ,
      layer4_out_conc_207_0})) * $signed((w5_rsci_idat[119:115]));
  assign Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_131_nl = conv_s2s_11_16(readslicef_15_11_4(Product1_1_124_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_125_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_116_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_117_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_120_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_121_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_112_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_113_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_110_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_111_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_12_16({Accum2_1_acc_390_nl , (Product1_1_107_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_itm_14_4_1[5:0])})
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_108_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_109_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_126_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_105_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_106_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_127_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_128_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_122_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_123_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_118_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_119_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_114_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_115_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));
  assign Accum2_1_acc_131_nl = nl_Accum2_1_acc_131_nl[15:0];
  assign nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_217_9 , layer4_out_conc_217_8_1 ,
      layer4_out_conc_217_0})) * $signed((w5_rsci_idat[194:190]));
  assign Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_219_9 , layer4_out_conc_219_8_1 ,
      layer4_out_conc_219_0})) * $signed((w5_rsci_idat[209:205]));
  assign Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_209_9 , layer4_out_conc_209_8_1 ,
      layer4_out_conc_209_0})) * $signed((w5_rsci_idat[134:130]));
  assign Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_211_9 , layer4_out_conc_211_8_1 ,
      layer4_out_conc_211_0})) * $signed((w5_rsci_idat[149:145]));
  assign Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_233_9 , layer4_out_conc_233_8_1 ,
      layer4_out_conc_233_0})) * $signed((w5_rsci_idat[314:310]));
  assign Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_235_9 , layer4_out_conc_235_8_1 ,
      layer4_out_conc_235_0})) * $signed((w5_rsci_idat[329:325]));
  assign Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_225_9 , layer4_out_conc_225_8_1 ,
      layer4_out_conc_225_0})) * $signed((w5_rsci_idat[254:250]));
  assign Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_227_9 , layer4_out_conc_227_8_1 ,
      layer4_out_conc_227_0})) * $signed((w5_rsci_idat[269:265]));
  assign Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_229_9 , layer4_out_conc_229_8_1 ,
      layer4_out_conc_229_0})) * $signed((w5_rsci_idat[284:280]));
  assign Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_231_9 , layer4_out_conc_231_8_1 ,
      layer4_out_conc_231_0})) * $signed((w5_rsci_idat[299:295]));
  assign Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_241_9 , layer4_out_conc_241_8_1 ,
      layer4_out_conc_241_0})) * $signed((w5_rsci_idat[374:370]));
  assign Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_243_9 , layer4_out_conc_243_8_1 ,
      layer4_out_conc_243_0})) * $signed((w5_rsci_idat[389:385]));
  assign Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_245_9 , layer4_out_conc_245_8_1 ,
      layer4_out_conc_245_0})) * $signed((w5_rsci_idat[404:400]));
  assign Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_247_9 , layer4_out_conc_247_8_1 ,
      layer4_out_conc_247_0})) * $signed((w5_rsci_idat[419:415]));
  assign Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_249_9 , layer4_out_conc_249_8_1 ,
      layer4_out_conc_249_0})) * $signed((w5_rsci_idat[434:430]));
  assign Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_251_9 , layer4_out_conc_251_8_1 ,
      layer4_out_conc_251_0})) * $signed((w5_rsci_idat[449:445]));
  assign Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_253_9 , layer4_out_conc_253_8_1 ,
      layer4_out_conc_253_0})) * $signed((w5_rsci_idat[464:460]));
  assign Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_255_9 , layer4_out_conc_255_8_1 ,
      layer4_out_conc_255_0})) * $signed((w5_rsci_idat[479:475]));
  assign Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_265_9 , layer4_out_conc_265_8_1 ,
      layer4_out_conc_265_0})) * $signed((w5_rsci_idat[554:550]));
  assign Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_267_9 , layer4_out_conc_267_8_1 ,
      layer4_out_conc_267_0})) * $signed((w5_rsci_idat[569:565]));
  assign Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_269_9 , layer4_out_conc_269_8_1 ,
      layer4_out_conc_269_0})) * $signed((w5_rsci_idat[584:580]));
  assign Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_271_9 , layer4_out_conc_271_8_1 ,
      layer4_out_conc_271_0})) * $signed((w5_rsci_idat[599:595]));
  assign Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_257_9 , layer4_out_conc_257_8_1 ,
      layer4_out_conc_257_0})) * $signed((w5_rsci_idat[494:490]));
  assign Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_259_9 , layer4_out_conc_259_8_1 ,
      layer4_out_conc_259_0})) * $signed((w5_rsci_idat[509:505]));
  assign Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_261_9 , layer4_out_conc_261_8_1 ,
      layer4_out_conc_261_0})) * $signed((w5_rsci_idat[524:520]));
  assign Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_263_9 , layer4_out_conc_263_8_1 ,
      layer4_out_conc_263_0})) * $signed((w5_rsci_idat[539:535]));
  assign Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_213_9 , layer4_out_conc_213_8_1 ,
      layer4_out_conc_213_0})) * $signed((w5_rsci_idat[164:160]));
  assign Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_215_9 , layer4_out_conc_215_8_1 ,
      layer4_out_conc_215_0})) * $signed((w5_rsci_idat[179:175]));
  assign Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_221_9 , layer4_out_conc_221_8_1 ,
      layer4_out_conc_221_0})) * $signed((w5_rsci_idat[224:220]));
  assign Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_223_9 , layer4_out_conc_223_8_1 ,
      layer4_out_conc_223_0})) * $signed((w5_rsci_idat[239:235]));
  assign Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_237_9 , layer4_out_conc_237_8_1 ,
      layer4_out_conc_237_0})) * $signed((w5_rsci_idat[344:340]));
  assign Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_239_9 , layer4_out_conc_239_8_1 ,
      layer4_out_conc_239_0})) * $signed((w5_rsci_idat[359:355]));
  assign Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl[14:0];
  assign nl_layer6_out_rsci_idat_47_32  = Accum2_1_acc_132_nl + Accum2_1_acc_131_nl
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config5_weight_t_product_mul_nl));

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [10:0] readslicef_15_11_4;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_15_11_4 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [15:0] readslicef_20_16_4;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_20_16_4 = tmp[15:0];
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_5_10 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_10 = {{5{vector[4]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_11_16 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_16 = {{5{vector[10]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_12_16 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_16 = {{4{vector[11]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    myproject
// ------------------------------------------------------------------


module myproject (
  clk, rst, input_1_rsc_dat, layer6_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer6_out_rsc_dat;
  input [8959:0] w2_rsc_dat;
  input [639:0] b2_rsc_dat;
  input [1919:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  converterBlock_myproject_core myproject_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .layer6_out_rsc_dat(layer6_out_rsc_dat),
      .w2_rsc_dat(w2_rsc_dat),
      .b2_rsc_dat(b2_rsc_dat),
      .w5_rsc_dat(w5_rsc_dat),
      .b5_rsc_dat(b5_rsc_dat)
    );
endmodule



