
//------> ./myproject_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module converterBlock_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./myproject_ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module converterBlock_ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./myproject_ROM_1i11_1o5_4ed11b0fc67dff9823222c14315e503abd.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
//
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Mon Oct 24 20:34:30 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i11_1o5_4ed11b0fc67dff9823222c14315e503abd
// ------------------------------------------------------------------


module converterBlock_ROM_1i11_1o5_4ed11b0fc67dff9823222c14315e503abd (
  I_1, O_1
);
  input [10:0] I_1;
  output [4:0] O_1;



  // Interconnect Declarations for Component Instantiations
  assign O_1 = MUX_v_5_1792_2(5'b11110, 5'b11011, 5'b11100, 5'b00010, 5'b01000, 5'b11010,
      5'b11110, 5'b00110, 5'b00000, 5'b00001, 5'b00001, 5'b00000, 5'b11100, 5'b11110,
      5'b00111, 5'b00111, 5'b10000, 5'b00110, 5'b00000, 5'b10101, 5'b11100, 5'b01000,
      5'b00000, 5'b00100, 5'b00110, 5'b00000, 5'b00011, 5'b00001, 5'b00001, 5'b00110,
      5'b00101, 5'b10110, 5'b11010, 5'b00001, 5'b00011, 5'b00011, 5'b00001, 5'b00011,
      5'b00011, 5'b00001, 5'b11111, 5'b11100, 5'b00000, 5'b00001, 5'b00001, 5'b11110,
      5'b11011, 5'b11110, 5'b11100, 5'b10111, 5'b11111, 5'b00000, 5'b00011, 5'b11111,
      5'b11111, 5'b11111, 5'b00000, 5'b11110, 5'b00000, 5'b10101, 5'b11000, 5'b11111,
      5'b00010, 5'b11001, 5'b00000, 5'b00000, 5'b11110, 5'b00000, 5'b11010, 5'b00010,
      5'b01101, 5'b00000, 5'b11111, 5'b00000, 5'b11111, 5'b00001, 5'b00011, 5'b11101,
      5'b00001, 5'b00011, 5'b00010, 5'b00001, 5'b11110, 5'b00000, 5'b00001, 5'b10011,
      5'b11011, 5'b00001, 5'b00001, 5'b00100, 5'b00101, 5'b00000, 5'b00000, 5'b00000,
      5'b11101, 5'b11011, 5'b01110, 5'b00001, 5'b11111, 5'b11111, 5'b11111, 5'b00000,
      5'b11111, 5'b11111, 5'b00000, 5'b01101, 5'b11001, 5'b00100, 5'b11110, 5'b00000,
      5'b11100, 5'b11011, 5'b11010, 5'b00000, 5'b01000, 5'b00011, 5'b11010, 5'b00010,
      5'b00001, 5'b00101, 5'b01000, 5'b00001, 5'b00101, 5'b11111, 5'b11001, 5'b11100,
      5'b00000, 5'b00101, 5'b11000, 5'b10001, 5'b11111, 5'b00000, 5'b11111, 5'b00111,
      5'b00110, 5'b00110, 5'b11111, 5'b11110, 5'b11100, 5'b11111, 5'b00000, 5'b00110,
      5'b00000, 5'b11110, 5'b00001, 5'b11110, 5'b11110, 5'b11111, 5'b11100, 5'b11011,
      5'b00010, 5'b01011, 5'b00001, 5'b11111, 5'b00100, 5'b11111, 5'b11111, 5'b00000,
      5'b11100, 5'b00010, 5'b00010, 5'b01111, 5'b11111, 5'b00010, 5'b00000, 5'b00000,
      5'b11100, 5'b11111, 5'b01011, 5'b10011, 5'b00000, 5'b11110, 5'b00000, 5'b11110,
      5'b11111, 5'b11100, 5'b00011, 5'b01100, 5'b11111, 5'b00101, 5'b11101, 5'b11111,
      5'b01001, 5'b11111, 5'b00000, 5'b01100, 5'b00000, 5'b00100, 5'b01111, 5'b11111,
      5'b00100, 5'b01000, 5'b11111, 5'b00000, 5'b00011, 5'b11111, 5'b11100, 5'b10000,
      5'b11001, 5'b11100, 5'b11011, 5'b00000, 5'b11111, 5'b11110, 5'b00101, 5'b11110,
      5'b00010, 5'b00111, 5'b00100, 5'b11111, 5'b00011, 5'b00001, 5'b11110, 5'b11101,
      5'b11001, 5'b01100, 5'b11111, 5'b00000, 5'b00101, 5'b11110, 5'b11111, 5'b00110,
      5'b10110, 5'b00010, 5'b10000, 5'b00000, 5'b11110, 5'b01000, 5'b00001, 5'b11111,
      5'b00000, 5'b00010, 5'b11101, 5'b10000, 5'b11110, 5'b00110, 5'b11000, 5'b11101,
      5'b00000, 5'b00101, 5'b00000, 5'b11111, 5'b11111, 5'b11010, 5'b11110, 5'b11110,
      5'b11111, 5'b01010, 5'b00001, 5'b11111, 5'b11111, 5'b01111, 5'b01111, 5'b01010,
      5'b11011, 5'b00010, 5'b10000, 5'b00011, 5'b11110, 5'b11010, 5'b11101, 5'b00010,
      5'b00010, 5'b00001, 5'b00010, 5'b11111, 5'b11101, 5'b11001, 5'b00011, 5'b01001,
      5'b00011, 5'b00110, 5'b11001, 5'b00000, 5'b11111, 5'b00100, 5'b10100, 5'b11110,
      5'b11110, 5'b11101, 5'b11101, 5'b11110, 5'b11111, 5'b00101, 5'b00010, 5'b00000,
      5'b11001, 5'b01111, 5'b11110, 5'b00010, 5'b11111, 5'b01111, 5'b11111, 5'b00001,
      5'b00101, 5'b11100, 5'b00001, 5'b00010, 5'b00100, 5'b11111, 5'b00001, 5'b11100,
      5'b00001, 5'b11111, 5'b01111, 5'b11010, 5'b10000, 5'b11100, 5'b10000, 5'b01000,
      5'b01111, 5'b01010, 5'b11111, 5'b00010, 5'b10101, 5'b00010, 5'b00011, 5'b00010,
      5'b00001, 5'b01011, 5'b00001, 5'b11101, 5'b11111, 5'b00010, 5'b01000, 5'b01111,
      5'b10011, 5'b00000, 5'b10000, 5'b00010, 5'b00101, 5'b11111, 5'b01000, 5'b00001,
      5'b11100, 5'b00101, 5'b01011, 5'b11110, 5'b11110, 5'b00001, 5'b00011, 5'b01010,
      5'b00100, 5'b00000, 5'b00000, 5'b01110, 5'b00011, 5'b00101, 5'b00000, 5'b01010,
      5'b01111, 5'b00011, 5'b01101, 5'b11001, 5'b00010, 5'b10111, 5'b10010, 5'b00001,
      5'b00010, 5'b11101, 5'b01110, 5'b01100, 5'b00100, 5'b00010, 5'b01000, 5'b00101,
      5'b10101, 5'b00011, 5'b10110, 5'b00100, 5'b11110, 5'b11100, 5'b00100, 5'b11111,
      5'b11110, 5'b11110, 5'b00011, 5'b00001, 5'b11010, 5'b00101, 5'b00000, 5'b00001,
      5'b00001, 5'b11100, 5'b01111, 5'b11000, 5'b10111, 5'b10000, 5'b01111, 5'b11101,
      5'b11100, 5'b00101, 5'b01111, 5'b11110, 5'b10100, 5'b11000, 5'b11101, 5'b11100,
      5'b10010, 5'b00100, 5'b01111, 5'b00101, 5'b11101, 5'b01111, 5'b11100, 5'b10100,
      5'b11000, 5'b11011, 5'b00000, 5'b00100, 5'b11001, 5'b10000, 5'b10001, 5'b00001,
      5'b10110, 5'b00111, 5'b00011, 5'b00010, 5'b00011, 5'b01010, 5'b11100, 5'b01111,
      5'b11000, 5'b01100, 5'b00001, 5'b10100, 5'b00010, 5'b01001, 5'b01111, 5'b10110,
      5'b00111, 5'b10110, 5'b00110, 5'b01001, 5'b00001, 5'b10100, 5'b11110, 5'b11001,
      5'b11101, 5'b10111, 5'b00001, 5'b01100, 5'b10101, 5'b00101, 5'b10000, 5'b00001,
      5'b11101, 5'b00111, 5'b11111, 5'b11110, 5'b11101, 5'b00100, 5'b00001, 5'b11111,
      5'b00010, 5'b11010, 5'b00010, 5'b00101, 5'b00100, 5'b11000, 5'b11101, 5'b01110,
      5'b00011, 5'b00001, 5'b00000, 5'b00110, 5'b11010, 5'b10000, 5'b11110, 5'b01111,
      5'b10001, 5'b00011, 5'b00100, 5'b00000, 5'b00110, 5'b00000, 5'b00011, 5'b11111,
      5'b11111, 5'b00011, 5'b11000, 5'b11011, 5'b10110, 5'b10001, 5'b00100, 5'b00110,
      5'b00101, 5'b00000, 5'b11010, 5'b00001, 5'b11111, 5'b01010, 5'b00000, 5'b00111,
      5'b11100, 5'b11010, 5'b10101, 5'b11001, 5'b10000, 5'b01000, 5'b10000, 5'b11010,
      5'b00000, 5'b00111, 5'b01001, 5'b00110, 5'b10100, 5'b01001, 5'b00100, 5'b11101,
      5'b11111, 5'b11100, 5'b11100, 5'b01111, 5'b00001, 5'b00001, 5'b01110, 5'b11011,
      5'b10000, 5'b11100, 5'b10111, 5'b01010, 5'b11000, 5'b10001, 5'b00000, 5'b10110,
      5'b11001, 5'b11110, 5'b00101, 5'b00000, 5'b01001, 5'b10000, 5'b01001, 5'b01111,
      5'b11000, 5'b11111, 5'b00011, 5'b00001, 5'b10101, 5'b10000, 5'b00000, 5'b01011,
      5'b11110, 5'b00010, 5'b00101, 5'b11110, 5'b00010, 5'b00000, 5'b01110, 5'b01111,
      5'b01010, 5'b11011, 5'b00010, 5'b01111, 5'b00100, 5'b10000, 5'b11010, 5'b00000,
      5'b01000, 5'b10111, 5'b11010, 5'b11100, 5'b11110, 5'b11001, 5'b00010, 5'b10000,
      5'b00101, 5'b11101, 5'b11000, 5'b00110, 5'b00000, 5'b01011, 5'b10101, 5'b00100,
      5'b11000, 5'b10111, 5'b00101, 5'b01101, 5'b10110, 5'b10101, 5'b11011, 5'b10101,
      5'b00111, 5'b10100, 5'b10011, 5'b00111, 5'b11110, 5'b11101, 5'b11011, 5'b10000,
      5'b00100, 5'b00001, 5'b00010, 5'b11110, 5'b01010, 5'b11100, 5'b10000, 5'b00110,
      5'b11010, 5'b00001, 5'b00000, 5'b00011, 5'b11101, 5'b00011, 5'b01111, 5'b00001,
      5'b10000, 5'b11101, 5'b00010, 5'b11100, 5'b01001, 5'b11000, 5'b01101, 5'b10000,
      5'b11011, 5'b11110, 5'b10011, 5'b11100, 5'b00101, 5'b00000, 5'b00010, 5'b00100,
      5'b00010, 5'b10000, 5'b11100, 5'b00001, 5'b11101, 5'b11110, 5'b10110, 5'b01100,
      5'b01011, 5'b10111, 5'b00101, 5'b11001, 5'b10100, 5'b00000, 5'b00110, 5'b10000,
      5'b11010, 5'b00101, 5'b00100, 5'b00000, 5'b01111, 5'b11111, 5'b10001, 5'b11111,
      5'b10011, 5'b10000, 5'b11010, 5'b00010, 5'b11010, 5'b00110, 5'b11101, 5'b00010,
      5'b01011, 5'b11101, 5'b11010, 5'b00011, 5'b11110, 5'b11011, 5'b01111, 5'b10100,
      5'b11001, 5'b11111, 5'b11101, 5'b00100, 5'b10100, 5'b01011, 5'b01110, 5'b10010,
      5'b10110, 5'b00101, 5'b11100, 5'b00100, 5'b00110, 5'b11011, 5'b11110, 5'b10101,
      5'b11010, 5'b11011, 5'b00001, 5'b01111, 5'b00100, 5'b10111, 5'b11111, 5'b10111,
      5'b11011, 5'b01111, 5'b10001, 5'b00100, 5'b11010, 5'b00011, 5'b11011, 5'b11101,
      5'b00001, 5'b11101, 5'b11111, 5'b00100, 5'b00001, 5'b10110, 5'b11011, 5'b00001,
      5'b11010, 5'b01001, 5'b00100, 5'b00010, 5'b11001, 5'b01100, 5'b11101, 5'b11011,
      5'b11100, 5'b11110, 5'b01010, 5'b11110, 5'b11010, 5'b01111, 5'b00000, 5'b11011,
      5'b00010, 5'b00000, 5'b00000, 5'b01010, 5'b00010, 5'b00010, 5'b01000, 5'b10101,
      5'b11101, 5'b00010, 5'b00100, 5'b00001, 5'b10000, 5'b00011, 5'b10000, 5'b11110,
      5'b00000, 5'b00010, 5'b10000, 5'b11000, 5'b00111, 5'b10000, 5'b10000, 5'b11110,
      5'b10000, 5'b11010, 5'b11011, 5'b01111, 5'b11101, 5'b10000, 5'b00001, 5'b10000,
      5'b00010, 5'b01111, 5'b00001, 5'b01111, 5'b11100, 5'b11101, 5'b01000, 5'b11010,
      5'b11110, 5'b10001, 5'b01000, 5'b01001, 5'b00001, 5'b00011, 5'b10000, 5'b11111,
      5'b11000, 5'b00011, 5'b01101, 5'b11010, 5'b11001, 5'b11100, 5'b10011, 5'b11101,
      5'b00010, 5'b01101, 5'b11000, 5'b11010, 5'b01111, 5'b01011, 5'b11101, 5'b11111,
      5'b11011, 5'b00000, 5'b10001, 5'b11100, 5'b11100, 5'b10000, 5'b10000, 5'b00000,
      5'b01111, 5'b10110, 5'b10011, 5'b00001, 5'b10110, 5'b01000, 5'b01011, 5'b10000,
      5'b01111, 5'b00001, 5'b00100, 5'b11111, 5'b11010, 5'b10110, 5'b11101, 5'b00001,
      5'b00101, 5'b10011, 5'b00101, 5'b10000, 5'b00101, 5'b01100, 5'b11111, 5'b10111,
      5'b10000, 5'b10001, 5'b00011, 5'b11010, 5'b00011, 5'b00110, 5'b11111, 5'b00100,
      5'b00011, 5'b11001, 5'b11000, 5'b10000, 5'b00011, 5'b10000, 5'b00101, 5'b00100,
      5'b11100, 5'b11011, 5'b00001, 5'b10011, 5'b10111, 5'b11000, 5'b10101, 5'b01100,
      5'b00101, 5'b01111, 5'b11011, 5'b10000, 5'b10000, 5'b10111, 5'b10111, 5'b00111,
      5'b00101, 5'b00100, 5'b00100, 5'b10101, 5'b00110, 5'b01111, 5'b01000, 5'b10000,
      5'b01111, 5'b00010, 5'b00001, 5'b00001, 5'b01111, 5'b11111, 5'b10000, 5'b01000,
      5'b01110, 5'b01000, 5'b00010, 5'b11011, 5'b10000, 5'b01111, 5'b01010, 5'b01011,
      5'b11111, 5'b00010, 5'b11011, 5'b00000, 5'b00000, 5'b01101, 5'b00011, 5'b10000,
      5'b11110, 5'b11101, 5'b01111, 5'b10110, 5'b11100, 5'b10101, 5'b01000, 5'b10111,
      5'b10011, 5'b01100, 5'b10000, 5'b11110, 5'b11111, 5'b00101, 5'b11111, 5'b00110,
      5'b00011, 5'b00011, 5'b10111, 5'b00101, 5'b11011, 5'b00000, 5'b10011, 5'b00000,
      5'b01000, 5'b00010, 5'b10100, 5'b11101, 5'b01110, 5'b11010, 5'b11111, 5'b11110,
      5'b10000, 5'b11100, 5'b10010, 5'b11000, 5'b11000, 5'b01111, 5'b11101, 5'b00010,
      5'b01111, 5'b01010, 5'b00101, 5'b00001, 5'b01000, 5'b00101, 5'b10101, 5'b00000,
      5'b01111, 5'b00101, 5'b11010, 5'b11111, 5'b00010, 5'b00101, 5'b11001, 5'b11010,
      5'b00000, 5'b01011, 5'b10011, 5'b11100, 5'b00100, 5'b00000, 5'b11010, 5'b01001,
      5'b00000, 5'b00000, 5'b11110, 5'b00111, 5'b10000, 5'b11101, 5'b00000, 5'b00111,
      5'b00000, 5'b00010, 5'b10000, 5'b00001, 5'b00000, 5'b00110, 5'b01111, 5'b11111,
      5'b11101, 5'b00010, 5'b11111, 5'b11100, 5'b11001, 5'b00001, 5'b00111, 5'b11101,
      5'b00110, 5'b11110, 5'b11110, 5'b00010, 5'b11110, 5'b11101, 5'b11101, 5'b11111,
      5'b11111, 5'b11100, 5'b10101, 5'b00010, 5'b11101, 5'b00110, 5'b00100, 5'b11001,
      5'b00100, 5'b11111, 5'b00011, 5'b00100, 5'b11101, 5'b00101, 5'b00110, 5'b10000,
      5'b00100, 5'b00010, 5'b10111, 5'b11110, 5'b10011, 5'b01111, 5'b11111, 5'b00010,
      5'b00110, 5'b11100, 5'b01111, 5'b11111, 5'b00011, 5'b11111, 5'b00010, 5'b00110,
      5'b01011, 5'b00001, 5'b11100, 5'b00000, 5'b01001, 5'b00000, 5'b01000, 5'b10100,
      5'b10011, 5'b00100, 5'b10100, 5'b00001, 5'b11111, 5'b00000, 5'b00010, 5'b00010,
      5'b10100, 5'b00001, 5'b01111, 5'b01111, 5'b11010, 5'b11011, 5'b11100, 5'b00100,
      5'b00100, 5'b01011, 5'b11011, 5'b11000, 5'b11111, 5'b00000, 5'b00001, 5'b10010,
      5'b01000, 5'b11110, 5'b00110, 5'b00001, 5'b11101, 5'b00001, 5'b00000, 5'b11011,
      5'b11101, 5'b01111, 5'b11101, 5'b00111, 5'b00000, 5'b11111, 5'b11101, 5'b00000,
      5'b11011, 5'b10010, 5'b00010, 5'b11111, 5'b00000, 5'b00010, 5'b01001, 5'b11000,
      5'b01011, 5'b11110, 5'b11010, 5'b11100, 5'b00001, 5'b00000, 5'b11010, 5'b00101,
      5'b00001, 5'b11111, 5'b00011, 5'b10000, 5'b01101, 5'b11111, 5'b00100, 5'b00000,
      5'b10001, 5'b01111, 5'b11111, 5'b01111, 5'b11110, 5'b00000, 5'b00000, 5'b01111,
      5'b00010, 5'b00000, 5'b00000, 5'b11011, 5'b00000, 5'b00100, 5'b00011, 5'b11111,
      5'b10110, 5'b11110, 5'b11000, 5'b00001, 5'b00100, 5'b00000, 5'b11110, 5'b11000,
      5'b01111, 5'b10111, 5'b11000, 5'b00000, 5'b11110, 5'b00001, 5'b11111, 5'b11111,
      5'b11011, 5'b11111, 5'b11001, 5'b00000, 5'b01010, 5'b11110, 5'b00001, 5'b01111,
      5'b10000, 5'b00101, 5'b00000, 5'b00001, 5'b11100, 5'b00000, 5'b11011, 5'b11001,
      5'b11110, 5'b00010, 5'b11110, 5'b10000, 5'b11001, 5'b00001, 5'b00000, 5'b00011,
      5'b00101, 5'b11111, 5'b11111, 5'b10000, 5'b00000, 5'b00001, 5'b00001, 5'b00100,
      5'b11110, 5'b11111, 5'b00100, 5'b00001, 5'b00000, 5'b10000, 5'b11110, 5'b11111,
      5'b11011, 5'b00001, 5'b10000, 5'b01000, 5'b00000, 5'b11111, 5'b00001, 5'b01011,
      5'b11111, 5'b10010, 5'b10110, 5'b00000, 5'b00001, 5'b01000, 5'b11010, 5'b11101,
      5'b00110, 5'b01000, 5'b10011, 5'b00100, 5'b00111, 5'b11111, 5'b00000, 5'b11100,
      5'b00000, 5'b00110, 5'b00010, 5'b00011, 5'b11110, 5'b11111, 5'b11010, 5'b00000,
      5'b11101, 5'b10111, 5'b00101, 5'b00001, 5'b11111, 5'b00110, 5'b11110, 5'b00010,
      5'b11011, 5'b00110, 5'b00001, 5'b01101, 5'b00000, 5'b11111, 5'b00011, 5'b00000,
      5'b11001, 5'b11001, 5'b11111, 5'b00100, 5'b11000, 5'b11110, 5'b11110, 5'b11111,
      5'b01111, 5'b11001, 5'b00011, 5'b10100, 5'b00000, 5'b00000, 5'b11111, 5'b00111,
      5'b11110, 5'b01110, 5'b11111, 5'b00001, 5'b11111, 5'b01011, 5'b10011, 5'b00001,
      5'b01111, 5'b00001, 5'b11101, 5'b01111, 5'b11110, 5'b11001, 5'b00111, 5'b01111,
      5'b10000, 5'b00001, 5'b00000, 5'b11111, 5'b11111, 5'b11111, 5'b11100, 5'b00101,
      5'b00110, 5'b00001, 5'b11101, 5'b11111, 5'b00010, 5'b00000, 5'b00000, 5'b10100,
      5'b10000, 5'b11101, 5'b11001, 5'b11100, 5'b11111, 5'b10000, 5'b11111, 5'b00111,
      5'b11111, 5'b00100, 5'b00000, 5'b10110, 5'b00010, 5'b10101, 5'b00000, 5'b11100,
      5'b11111, 5'b11100, 5'b11010, 5'b11100, 5'b11111, 5'b11011, 5'b00011, 5'b10000,
      5'b00000, 5'b01000, 5'b11111, 5'b01111, 5'b00000, 5'b00000, 5'b11100, 5'b11111,
      5'b00000, 5'b00101, 5'b01111, 5'b10110, 5'b01101, 5'b00000, 5'b10100, 5'b11010,
      5'b00110, 5'b00001, 5'b00011, 5'b00000, 5'b01101, 5'b11010, 5'b11100, 5'b00010,
      5'b11000, 5'b00001, 5'b11101, 5'b00011, 5'b11101, 5'b00000, 5'b11110, 5'b10101,
      5'b10010, 5'b00001, 5'b11101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000,
      5'b01111, 5'b00110, 5'b00010, 5'b00000, 5'b00000, 5'b10011, 5'b11100, 5'b01000,
      5'b11100, 5'b00011, 5'b00010, 5'b11001, 5'b11110, 5'b00000, 5'b01101, 5'b01000,
      5'b00010, 5'b00100, 5'b11001, 5'b11111, 5'b00000, 5'b00010, 5'b00000, 5'b00000,
      5'b11110, 5'b00000, 5'b11101, 5'b11101, 5'b00001, 5'b00000, 5'b00000, 5'b00000,
      5'b00000, 5'b10010, 5'b11100, 5'b11111, 5'b00001, 5'b11011, 5'b01100, 5'b11111,
      5'b11110, 5'b11101, 5'b01001, 5'b10101, 5'b00010, 5'b00101, 5'b10110, 5'b11011,
      5'b01011, 5'b00100, 5'b00010, 5'b00000, 5'b11111, 5'b00000, 5'b01111, 5'b01110,
      5'b00111, 5'b00000, 5'b11101, 5'b11111, 5'b01001, 5'b11111, 5'b00000, 5'b11010,
      5'b01111, 5'b11111, 5'b00010, 5'b00011, 5'b00010, 5'b11011, 5'b00001, 5'b00001,
      5'b11110, 5'b00100, 5'b00111, 5'b01001, 5'b11111, 5'b01101, 5'b11111, 5'b01010,
      5'b01000, 5'b00001, 5'b11101, 5'b01011, 5'b00110, 5'b00000, 5'b11011, 5'b01001,
      5'b00010, 5'b00011, 5'b00010, 5'b10000, 5'b11111, 5'b11110, 5'b10110, 5'b00000,
      5'b11111, 5'b00100, 5'b11101, 5'b01101, 5'b10001, 5'b00000, 5'b10101, 5'b11011,
      5'b10010, 5'b01001, 5'b00000, 5'b00001, 5'b00100, 5'b01000, 5'b11100, 5'b11101,
      5'b00000, 5'b00111, 5'b01000, 5'b00011, 5'b00010, 5'b01000, 5'b00111, 5'b01010,
      5'b11111, 5'b11111, 5'b11101, 5'b00011, 5'b00001, 5'b00000, 5'b00010, 5'b11111,
      5'b00001, 5'b00001, 5'b00100, 5'b11111, 5'b00000, 5'b01010, 5'b00011, 5'b10111,
      5'b00000, 5'b11000, 5'b11110, 5'b11111, 5'b11110, 5'b11111, 5'b10000, 5'b11101,
      5'b00001, 5'b00000, 5'b11010, 5'b00000, 5'b00000, 5'b11101, 5'b00101, 5'b11110,
      5'b00100, 5'b11111, 5'b01010, 5'b11110, 5'b00001, 5'b01100, 5'b10010, 5'b11110,
      5'b00000, 5'b00111, 5'b11111, 5'b11011, 5'b11011, 5'b00110, 5'b10101, 5'b01100,
      5'b10001, 5'b00000, 5'b11111, 5'b00011, 5'b11101, 5'b11100, 5'b00111, 5'b11111,
      5'b01111, 5'b00011, 5'b11110, 5'b11111, 5'b00011, 5'b11110, 5'b11010, 5'b01001,
      5'b11101, 5'b00011, 5'b00011, 5'b11110, 5'b11111, 5'b00110, 5'b00000, 5'b00100,
      5'b00101, 5'b11110, 5'b11100, 5'b00000, 5'b11110, 5'b11101, 5'b11001, 5'b10111,
      5'b11111, 5'b11110, 5'b00110, 5'b11101, 5'b00010, 5'b11010, 5'b00101, 5'b00101,
      5'b00100, 5'b00000, 5'b01111, 5'b00000, 5'b11011, 5'b11111, 5'b11001, 5'b11011,
      5'b00010, 5'b00001, 5'b10100, 5'b00110, 5'b00000, 5'b11111, 5'b01111, 5'b00000,
      5'b00010, 5'b11101, 5'b10100, 5'b10100, 5'b00000, 5'b00000, 5'b00101, 5'b11010,
      5'b11111, 5'b00011, 5'b11111, 5'b11111, 5'b11111, 5'b11010, 5'b11110, 5'b00000,
      5'b11111, 5'b00000, 5'b00101, 5'b00110, 5'b00010, 5'b00001, 5'b11011, 5'b11100,
      5'b11100, 5'b11110, 5'b00101, 5'b11100, 5'b11010, 5'b00000, 5'b11110, 5'b00000,
      5'b10100, 5'b11101, 5'b11100, 5'b11001, 5'b11110, 5'b00001, 5'b00101, 5'b00010,
      5'b00000, 5'b11110, 5'b11001, 5'b11100, 5'b00100, 5'b11111, 5'b01010, 5'b00010,
      5'b11000, 5'b11111, 5'b01010, 5'b10110, 5'b00000, 5'b00010, 5'b11000, 5'b00000,
      5'b00000, 5'b00110, 5'b11101, 5'b01111, 5'b00001, 5'b10111, 5'b01100, 5'b11111,
      5'b00001, 5'b11011, 5'b00101, 5'b00100, 5'b00011, 5'b11110, 5'b00100, 5'b00010,
      5'b00100, 5'b00000, 5'b11111, 5'b11101, 5'b00000, 5'b00001, 5'b11101, 5'b11010,
      5'b11000, 5'b00001, 5'b10111, 5'b00110, 5'b11111, 5'b11001, 5'b00100, 5'b00010,
      5'b00000, 5'b11111, 5'b00010, 5'b00000, 5'b11101, 5'b00000, 5'b11111, 5'b00001,
      5'b10110, 5'b00000, 5'b00001, 5'b11101, 5'b00001, 5'b00100, 5'b00010, 5'b00000,
      5'b00001, 5'b00100, 5'b00000, 5'b11010, 5'b00111, 5'b11001, 5'b00001, 5'b11101,
      5'b00010, 5'b11110, 5'b01011, 5'b11001, 5'b11111, 5'b00100, 5'b00101, 5'b00101,
      5'b11111, 5'b00000, 5'b00011, 5'b11111, 5'b00000, 5'b00100, 5'b00001, 5'b00000,
      5'b00101, 5'b00010, 5'b01001, 5'b01001, 5'b11110, 5'b11110, 5'b10111, 5'b11100,
      5'b00011, 5'b01000, 5'b10111, 5'b10001, 5'b11011, 5'b11100, 5'b00001, 5'b10110,
      5'b00011, 5'b11100, 5'b10101, 5'b11101, 5'b11000, 5'b10110, 5'b00111, 5'b11111,
      5'b11010, 5'b11011, 5'b10000, 5'b10111, 5'b11111, 5'b01000, 5'b11110, 5'b00001,
      5'b10011, 5'b00001, 5'b00010, 5'b01111, 5'b00001, 5'b01101, 5'b01011, 5'b11110,
      5'b01111, 5'b10000, 5'b11100, 5'b10100, 5'b00010, 5'b00011, 5'b10001, 5'b11000,
      5'b00100, 5'b10111, 5'b00101, 5'b00110, 5'b11101, 5'b10110, 5'b01111, 5'b00101,
      5'b00111, 5'b11001, 5'b00001, 5'b01011, 5'b10111, 5'b01000, 5'b10111, 5'b01111,
      5'b00101, 5'b01111, 5'b10011, 5'b11000, 5'b11101, 5'b01111, 5'b11000, 5'b10000,
      5'b01011, 5'b11010, 5'b11000, 5'b00100, 5'b00011, 5'b10001, 5'b11001, 5'b00001,
      5'b00011, 5'b00111, 5'b00101, 5'b10101, 5'b10010, 5'b01011, 5'b01001, 5'b11010,
      5'b11000, 5'b01100, 5'b00100, 5'b11001, 5'b00101, 5'b01111, 5'b00110, 5'b01110,
      5'b01011, 5'b11010, 5'b10000, 5'b00100, 5'b11011, 5'b10111, 5'b11111, 5'b00101,
      5'b00010, 5'b11100, 5'b11000, 5'b01001, 5'b00011, 5'b11101, 5'b11000, 5'b01011,
      5'b11111, 5'b11111, 5'b10100, 5'b01111, 5'b00101, 5'b00000, 5'b01001, 5'b10000,
      5'b11100, 5'b01110, 5'b01001, 5'b01111, 5'b11110, 5'b01110, 5'b00011, 5'b00001,
      5'b00001, 5'b00111, I_1);

  function automatic [4:0] MUX_v_5_1792_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [4:0] input_4;
    input [4:0] input_5;
    input [4:0] input_6;
    input [4:0] input_7;
    input [4:0] input_8;
    input [4:0] input_9;
    input [4:0] input_10;
    input [4:0] input_11;
    input [4:0] input_12;
    input [4:0] input_13;
    input [4:0] input_14;
    input [4:0] input_15;
    input [4:0] input_16;
    input [4:0] input_17;
    input [4:0] input_18;
    input [4:0] input_19;
    input [4:0] input_20;
    input [4:0] input_21;
    input [4:0] input_22;
    input [4:0] input_23;
    input [4:0] input_24;
    input [4:0] input_25;
    input [4:0] input_26;
    input [4:0] input_27;
    input [4:0] input_28;
    input [4:0] input_29;
    input [4:0] input_30;
    input [4:0] input_31;
    input [4:0] input_32;
    input [4:0] input_33;
    input [4:0] input_34;
    input [4:0] input_35;
    input [4:0] input_36;
    input [4:0] input_37;
    input [4:0] input_38;
    input [4:0] input_39;
    input [4:0] input_40;
    input [4:0] input_41;
    input [4:0] input_42;
    input [4:0] input_43;
    input [4:0] input_44;
    input [4:0] input_45;
    input [4:0] input_46;
    input [4:0] input_47;
    input [4:0] input_48;
    input [4:0] input_49;
    input [4:0] input_50;
    input [4:0] input_51;
    input [4:0] input_52;
    input [4:0] input_53;
    input [4:0] input_54;
    input [4:0] input_55;
    input [4:0] input_56;
    input [4:0] input_57;
    input [4:0] input_58;
    input [4:0] input_59;
    input [4:0] input_60;
    input [4:0] input_61;
    input [4:0] input_62;
    input [4:0] input_63;
    input [4:0] input_64;
    input [4:0] input_65;
    input [4:0] input_66;
    input [4:0] input_67;
    input [4:0] input_68;
    input [4:0] input_69;
    input [4:0] input_70;
    input [4:0] input_71;
    input [4:0] input_72;
    input [4:0] input_73;
    input [4:0] input_74;
    input [4:0] input_75;
    input [4:0] input_76;
    input [4:0] input_77;
    input [4:0] input_78;
    input [4:0] input_79;
    input [4:0] input_80;
    input [4:0] input_81;
    input [4:0] input_82;
    input [4:0] input_83;
    input [4:0] input_84;
    input [4:0] input_85;
    input [4:0] input_86;
    input [4:0] input_87;
    input [4:0] input_88;
    input [4:0] input_89;
    input [4:0] input_90;
    input [4:0] input_91;
    input [4:0] input_92;
    input [4:0] input_93;
    input [4:0] input_94;
    input [4:0] input_95;
    input [4:0] input_96;
    input [4:0] input_97;
    input [4:0] input_98;
    input [4:0] input_99;
    input [4:0] input_100;
    input [4:0] input_101;
    input [4:0] input_102;
    input [4:0] input_103;
    input [4:0] input_104;
    input [4:0] input_105;
    input [4:0] input_106;
    input [4:0] input_107;
    input [4:0] input_108;
    input [4:0] input_109;
    input [4:0] input_110;
    input [4:0] input_111;
    input [4:0] input_112;
    input [4:0] input_113;
    input [4:0] input_114;
    input [4:0] input_115;
    input [4:0] input_116;
    input [4:0] input_117;
    input [4:0] input_118;
    input [4:0] input_119;
    input [4:0] input_120;
    input [4:0] input_121;
    input [4:0] input_122;
    input [4:0] input_123;
    input [4:0] input_124;
    input [4:0] input_125;
    input [4:0] input_126;
    input [4:0] input_127;
    input [4:0] input_128;
    input [4:0] input_129;
    input [4:0] input_130;
    input [4:0] input_131;
    input [4:0] input_132;
    input [4:0] input_133;
    input [4:0] input_134;
    input [4:0] input_135;
    input [4:0] input_136;
    input [4:0] input_137;
    input [4:0] input_138;
    input [4:0] input_139;
    input [4:0] input_140;
    input [4:0] input_141;
    input [4:0] input_142;
    input [4:0] input_143;
    input [4:0] input_144;
    input [4:0] input_145;
    input [4:0] input_146;
    input [4:0] input_147;
    input [4:0] input_148;
    input [4:0] input_149;
    input [4:0] input_150;
    input [4:0] input_151;
    input [4:0] input_152;
    input [4:0] input_153;
    input [4:0] input_154;
    input [4:0] input_155;
    input [4:0] input_156;
    input [4:0] input_157;
    input [4:0] input_158;
    input [4:0] input_159;
    input [4:0] input_160;
    input [4:0] input_161;
    input [4:0] input_162;
    input [4:0] input_163;
    input [4:0] input_164;
    input [4:0] input_165;
    input [4:0] input_166;
    input [4:0] input_167;
    input [4:0] input_168;
    input [4:0] input_169;
    input [4:0] input_170;
    input [4:0] input_171;
    input [4:0] input_172;
    input [4:0] input_173;
    input [4:0] input_174;
    input [4:0] input_175;
    input [4:0] input_176;
    input [4:0] input_177;
    input [4:0] input_178;
    input [4:0] input_179;
    input [4:0] input_180;
    input [4:0] input_181;
    input [4:0] input_182;
    input [4:0] input_183;
    input [4:0] input_184;
    input [4:0] input_185;
    input [4:0] input_186;
    input [4:0] input_187;
    input [4:0] input_188;
    input [4:0] input_189;
    input [4:0] input_190;
    input [4:0] input_191;
    input [4:0] input_192;
    input [4:0] input_193;
    input [4:0] input_194;
    input [4:0] input_195;
    input [4:0] input_196;
    input [4:0] input_197;
    input [4:0] input_198;
    input [4:0] input_199;
    input [4:0] input_200;
    input [4:0] input_201;
    input [4:0] input_202;
    input [4:0] input_203;
    input [4:0] input_204;
    input [4:0] input_205;
    input [4:0] input_206;
    input [4:0] input_207;
    input [4:0] input_208;
    input [4:0] input_209;
    input [4:0] input_210;
    input [4:0] input_211;
    input [4:0] input_212;
    input [4:0] input_213;
    input [4:0] input_214;
    input [4:0] input_215;
    input [4:0] input_216;
    input [4:0] input_217;
    input [4:0] input_218;
    input [4:0] input_219;
    input [4:0] input_220;
    input [4:0] input_221;
    input [4:0] input_222;
    input [4:0] input_223;
    input [4:0] input_224;
    input [4:0] input_225;
    input [4:0] input_226;
    input [4:0] input_227;
    input [4:0] input_228;
    input [4:0] input_229;
    input [4:0] input_230;
    input [4:0] input_231;
    input [4:0] input_232;
    input [4:0] input_233;
    input [4:0] input_234;
    input [4:0] input_235;
    input [4:0] input_236;
    input [4:0] input_237;
    input [4:0] input_238;
    input [4:0] input_239;
    input [4:0] input_240;
    input [4:0] input_241;
    input [4:0] input_242;
    input [4:0] input_243;
    input [4:0] input_244;
    input [4:0] input_245;
    input [4:0] input_246;
    input [4:0] input_247;
    input [4:0] input_248;
    input [4:0] input_249;
    input [4:0] input_250;
    input [4:0] input_251;
    input [4:0] input_252;
    input [4:0] input_253;
    input [4:0] input_254;
    input [4:0] input_255;
    input [4:0] input_256;
    input [4:0] input_257;
    input [4:0] input_258;
    input [4:0] input_259;
    input [4:0] input_260;
    input [4:0] input_261;
    input [4:0] input_262;
    input [4:0] input_263;
    input [4:0] input_264;
    input [4:0] input_265;
    input [4:0] input_266;
    input [4:0] input_267;
    input [4:0] input_268;
    input [4:0] input_269;
    input [4:0] input_270;
    input [4:0] input_271;
    input [4:0] input_272;
    input [4:0] input_273;
    input [4:0] input_274;
    input [4:0] input_275;
    input [4:0] input_276;
    input [4:0] input_277;
    input [4:0] input_278;
    input [4:0] input_279;
    input [4:0] input_280;
    input [4:0] input_281;
    input [4:0] input_282;
    input [4:0] input_283;
    input [4:0] input_284;
    input [4:0] input_285;
    input [4:0] input_286;
    input [4:0] input_287;
    input [4:0] input_288;
    input [4:0] input_289;
    input [4:0] input_290;
    input [4:0] input_291;
    input [4:0] input_292;
    input [4:0] input_293;
    input [4:0] input_294;
    input [4:0] input_295;
    input [4:0] input_296;
    input [4:0] input_297;
    input [4:0] input_298;
    input [4:0] input_299;
    input [4:0] input_300;
    input [4:0] input_301;
    input [4:0] input_302;
    input [4:0] input_303;
    input [4:0] input_304;
    input [4:0] input_305;
    input [4:0] input_306;
    input [4:0] input_307;
    input [4:0] input_308;
    input [4:0] input_309;
    input [4:0] input_310;
    input [4:0] input_311;
    input [4:0] input_312;
    input [4:0] input_313;
    input [4:0] input_314;
    input [4:0] input_315;
    input [4:0] input_316;
    input [4:0] input_317;
    input [4:0] input_318;
    input [4:0] input_319;
    input [4:0] input_320;
    input [4:0] input_321;
    input [4:0] input_322;
    input [4:0] input_323;
    input [4:0] input_324;
    input [4:0] input_325;
    input [4:0] input_326;
    input [4:0] input_327;
    input [4:0] input_328;
    input [4:0] input_329;
    input [4:0] input_330;
    input [4:0] input_331;
    input [4:0] input_332;
    input [4:0] input_333;
    input [4:0] input_334;
    input [4:0] input_335;
    input [4:0] input_336;
    input [4:0] input_337;
    input [4:0] input_338;
    input [4:0] input_339;
    input [4:0] input_340;
    input [4:0] input_341;
    input [4:0] input_342;
    input [4:0] input_343;
    input [4:0] input_344;
    input [4:0] input_345;
    input [4:0] input_346;
    input [4:0] input_347;
    input [4:0] input_348;
    input [4:0] input_349;
    input [4:0] input_350;
    input [4:0] input_351;
    input [4:0] input_352;
    input [4:0] input_353;
    input [4:0] input_354;
    input [4:0] input_355;
    input [4:0] input_356;
    input [4:0] input_357;
    input [4:0] input_358;
    input [4:0] input_359;
    input [4:0] input_360;
    input [4:0] input_361;
    input [4:0] input_362;
    input [4:0] input_363;
    input [4:0] input_364;
    input [4:0] input_365;
    input [4:0] input_366;
    input [4:0] input_367;
    input [4:0] input_368;
    input [4:0] input_369;
    input [4:0] input_370;
    input [4:0] input_371;
    input [4:0] input_372;
    input [4:0] input_373;
    input [4:0] input_374;
    input [4:0] input_375;
    input [4:0] input_376;
    input [4:0] input_377;
    input [4:0] input_378;
    input [4:0] input_379;
    input [4:0] input_380;
    input [4:0] input_381;
    input [4:0] input_382;
    input [4:0] input_383;
    input [4:0] input_384;
    input [4:0] input_385;
    input [4:0] input_386;
    input [4:0] input_387;
    input [4:0] input_388;
    input [4:0] input_389;
    input [4:0] input_390;
    input [4:0] input_391;
    input [4:0] input_392;
    input [4:0] input_393;
    input [4:0] input_394;
    input [4:0] input_395;
    input [4:0] input_396;
    input [4:0] input_397;
    input [4:0] input_398;
    input [4:0] input_399;
    input [4:0] input_400;
    input [4:0] input_401;
    input [4:0] input_402;
    input [4:0] input_403;
    input [4:0] input_404;
    input [4:0] input_405;
    input [4:0] input_406;
    input [4:0] input_407;
    input [4:0] input_408;
    input [4:0] input_409;
    input [4:0] input_410;
    input [4:0] input_411;
    input [4:0] input_412;
    input [4:0] input_413;
    input [4:0] input_414;
    input [4:0] input_415;
    input [4:0] input_416;
    input [4:0] input_417;
    input [4:0] input_418;
    input [4:0] input_419;
    input [4:0] input_420;
    input [4:0] input_421;
    input [4:0] input_422;
    input [4:0] input_423;
    input [4:0] input_424;
    input [4:0] input_425;
    input [4:0] input_426;
    input [4:0] input_427;
    input [4:0] input_428;
    input [4:0] input_429;
    input [4:0] input_430;
    input [4:0] input_431;
    input [4:0] input_432;
    input [4:0] input_433;
    input [4:0] input_434;
    input [4:0] input_435;
    input [4:0] input_436;
    input [4:0] input_437;
    input [4:0] input_438;
    input [4:0] input_439;
    input [4:0] input_440;
    input [4:0] input_441;
    input [4:0] input_442;
    input [4:0] input_443;
    input [4:0] input_444;
    input [4:0] input_445;
    input [4:0] input_446;
    input [4:0] input_447;
    input [4:0] input_448;
    input [4:0] input_449;
    input [4:0] input_450;
    input [4:0] input_451;
    input [4:0] input_452;
    input [4:0] input_453;
    input [4:0] input_454;
    input [4:0] input_455;
    input [4:0] input_456;
    input [4:0] input_457;
    input [4:0] input_458;
    input [4:0] input_459;
    input [4:0] input_460;
    input [4:0] input_461;
    input [4:0] input_462;
    input [4:0] input_463;
    input [4:0] input_464;
    input [4:0] input_465;
    input [4:0] input_466;
    input [4:0] input_467;
    input [4:0] input_468;
    input [4:0] input_469;
    input [4:0] input_470;
    input [4:0] input_471;
    input [4:0] input_472;
    input [4:0] input_473;
    input [4:0] input_474;
    input [4:0] input_475;
    input [4:0] input_476;
    input [4:0] input_477;
    input [4:0] input_478;
    input [4:0] input_479;
    input [4:0] input_480;
    input [4:0] input_481;
    input [4:0] input_482;
    input [4:0] input_483;
    input [4:0] input_484;
    input [4:0] input_485;
    input [4:0] input_486;
    input [4:0] input_487;
    input [4:0] input_488;
    input [4:0] input_489;
    input [4:0] input_490;
    input [4:0] input_491;
    input [4:0] input_492;
    input [4:0] input_493;
    input [4:0] input_494;
    input [4:0] input_495;
    input [4:0] input_496;
    input [4:0] input_497;
    input [4:0] input_498;
    input [4:0] input_499;
    input [4:0] input_500;
    input [4:0] input_501;
    input [4:0] input_502;
    input [4:0] input_503;
    input [4:0] input_504;
    input [4:0] input_505;
    input [4:0] input_506;
    input [4:0] input_507;
    input [4:0] input_508;
    input [4:0] input_509;
    input [4:0] input_510;
    input [4:0] input_511;
    input [4:0] input_512;
    input [4:0] input_513;
    input [4:0] input_514;
    input [4:0] input_515;
    input [4:0] input_516;
    input [4:0] input_517;
    input [4:0] input_518;
    input [4:0] input_519;
    input [4:0] input_520;
    input [4:0] input_521;
    input [4:0] input_522;
    input [4:0] input_523;
    input [4:0] input_524;
    input [4:0] input_525;
    input [4:0] input_526;
    input [4:0] input_527;
    input [4:0] input_528;
    input [4:0] input_529;
    input [4:0] input_530;
    input [4:0] input_531;
    input [4:0] input_532;
    input [4:0] input_533;
    input [4:0] input_534;
    input [4:0] input_535;
    input [4:0] input_536;
    input [4:0] input_537;
    input [4:0] input_538;
    input [4:0] input_539;
    input [4:0] input_540;
    input [4:0] input_541;
    input [4:0] input_542;
    input [4:0] input_543;
    input [4:0] input_544;
    input [4:0] input_545;
    input [4:0] input_546;
    input [4:0] input_547;
    input [4:0] input_548;
    input [4:0] input_549;
    input [4:0] input_550;
    input [4:0] input_551;
    input [4:0] input_552;
    input [4:0] input_553;
    input [4:0] input_554;
    input [4:0] input_555;
    input [4:0] input_556;
    input [4:0] input_557;
    input [4:0] input_558;
    input [4:0] input_559;
    input [4:0] input_560;
    input [4:0] input_561;
    input [4:0] input_562;
    input [4:0] input_563;
    input [4:0] input_564;
    input [4:0] input_565;
    input [4:0] input_566;
    input [4:0] input_567;
    input [4:0] input_568;
    input [4:0] input_569;
    input [4:0] input_570;
    input [4:0] input_571;
    input [4:0] input_572;
    input [4:0] input_573;
    input [4:0] input_574;
    input [4:0] input_575;
    input [4:0] input_576;
    input [4:0] input_577;
    input [4:0] input_578;
    input [4:0] input_579;
    input [4:0] input_580;
    input [4:0] input_581;
    input [4:0] input_582;
    input [4:0] input_583;
    input [4:0] input_584;
    input [4:0] input_585;
    input [4:0] input_586;
    input [4:0] input_587;
    input [4:0] input_588;
    input [4:0] input_589;
    input [4:0] input_590;
    input [4:0] input_591;
    input [4:0] input_592;
    input [4:0] input_593;
    input [4:0] input_594;
    input [4:0] input_595;
    input [4:0] input_596;
    input [4:0] input_597;
    input [4:0] input_598;
    input [4:0] input_599;
    input [4:0] input_600;
    input [4:0] input_601;
    input [4:0] input_602;
    input [4:0] input_603;
    input [4:0] input_604;
    input [4:0] input_605;
    input [4:0] input_606;
    input [4:0] input_607;
    input [4:0] input_608;
    input [4:0] input_609;
    input [4:0] input_610;
    input [4:0] input_611;
    input [4:0] input_612;
    input [4:0] input_613;
    input [4:0] input_614;
    input [4:0] input_615;
    input [4:0] input_616;
    input [4:0] input_617;
    input [4:0] input_618;
    input [4:0] input_619;
    input [4:0] input_620;
    input [4:0] input_621;
    input [4:0] input_622;
    input [4:0] input_623;
    input [4:0] input_624;
    input [4:0] input_625;
    input [4:0] input_626;
    input [4:0] input_627;
    input [4:0] input_628;
    input [4:0] input_629;
    input [4:0] input_630;
    input [4:0] input_631;
    input [4:0] input_632;
    input [4:0] input_633;
    input [4:0] input_634;
    input [4:0] input_635;
    input [4:0] input_636;
    input [4:0] input_637;
    input [4:0] input_638;
    input [4:0] input_639;
    input [4:0] input_640;
    input [4:0] input_641;
    input [4:0] input_642;
    input [4:0] input_643;
    input [4:0] input_644;
    input [4:0] input_645;
    input [4:0] input_646;
    input [4:0] input_647;
    input [4:0] input_648;
    input [4:0] input_649;
    input [4:0] input_650;
    input [4:0] input_651;
    input [4:0] input_652;
    input [4:0] input_653;
    input [4:0] input_654;
    input [4:0] input_655;
    input [4:0] input_656;
    input [4:0] input_657;
    input [4:0] input_658;
    input [4:0] input_659;
    input [4:0] input_660;
    input [4:0] input_661;
    input [4:0] input_662;
    input [4:0] input_663;
    input [4:0] input_664;
    input [4:0] input_665;
    input [4:0] input_666;
    input [4:0] input_667;
    input [4:0] input_668;
    input [4:0] input_669;
    input [4:0] input_670;
    input [4:0] input_671;
    input [4:0] input_672;
    input [4:0] input_673;
    input [4:0] input_674;
    input [4:0] input_675;
    input [4:0] input_676;
    input [4:0] input_677;
    input [4:0] input_678;
    input [4:0] input_679;
    input [4:0] input_680;
    input [4:0] input_681;
    input [4:0] input_682;
    input [4:0] input_683;
    input [4:0] input_684;
    input [4:0] input_685;
    input [4:0] input_686;
    input [4:0] input_687;
    input [4:0] input_688;
    input [4:0] input_689;
    input [4:0] input_690;
    input [4:0] input_691;
    input [4:0] input_692;
    input [4:0] input_693;
    input [4:0] input_694;
    input [4:0] input_695;
    input [4:0] input_696;
    input [4:0] input_697;
    input [4:0] input_698;
    input [4:0] input_699;
    input [4:0] input_700;
    input [4:0] input_701;
    input [4:0] input_702;
    input [4:0] input_703;
    input [4:0] input_704;
    input [4:0] input_705;
    input [4:0] input_706;
    input [4:0] input_707;
    input [4:0] input_708;
    input [4:0] input_709;
    input [4:0] input_710;
    input [4:0] input_711;
    input [4:0] input_712;
    input [4:0] input_713;
    input [4:0] input_714;
    input [4:0] input_715;
    input [4:0] input_716;
    input [4:0] input_717;
    input [4:0] input_718;
    input [4:0] input_719;
    input [4:0] input_720;
    input [4:0] input_721;
    input [4:0] input_722;
    input [4:0] input_723;
    input [4:0] input_724;
    input [4:0] input_725;
    input [4:0] input_726;
    input [4:0] input_727;
    input [4:0] input_728;
    input [4:0] input_729;
    input [4:0] input_730;
    input [4:0] input_731;
    input [4:0] input_732;
    input [4:0] input_733;
    input [4:0] input_734;
    input [4:0] input_735;
    input [4:0] input_736;
    input [4:0] input_737;
    input [4:0] input_738;
    input [4:0] input_739;
    input [4:0] input_740;
    input [4:0] input_741;
    input [4:0] input_742;
    input [4:0] input_743;
    input [4:0] input_744;
    input [4:0] input_745;
    input [4:0] input_746;
    input [4:0] input_747;
    input [4:0] input_748;
    input [4:0] input_749;
    input [4:0] input_750;
    input [4:0] input_751;
    input [4:0] input_752;
    input [4:0] input_753;
    input [4:0] input_754;
    input [4:0] input_755;
    input [4:0] input_756;
    input [4:0] input_757;
    input [4:0] input_758;
    input [4:0] input_759;
    input [4:0] input_760;
    input [4:0] input_761;
    input [4:0] input_762;
    input [4:0] input_763;
    input [4:0] input_764;
    input [4:0] input_765;
    input [4:0] input_766;
    input [4:0] input_767;
    input [4:0] input_768;
    input [4:0] input_769;
    input [4:0] input_770;
    input [4:0] input_771;
    input [4:0] input_772;
    input [4:0] input_773;
    input [4:0] input_774;
    input [4:0] input_775;
    input [4:0] input_776;
    input [4:0] input_777;
    input [4:0] input_778;
    input [4:0] input_779;
    input [4:0] input_780;
    input [4:0] input_781;
    input [4:0] input_782;
    input [4:0] input_783;
    input [4:0] input_784;
    input [4:0] input_785;
    input [4:0] input_786;
    input [4:0] input_787;
    input [4:0] input_788;
    input [4:0] input_789;
    input [4:0] input_790;
    input [4:0] input_791;
    input [4:0] input_792;
    input [4:0] input_793;
    input [4:0] input_794;
    input [4:0] input_795;
    input [4:0] input_796;
    input [4:0] input_797;
    input [4:0] input_798;
    input [4:0] input_799;
    input [4:0] input_800;
    input [4:0] input_801;
    input [4:0] input_802;
    input [4:0] input_803;
    input [4:0] input_804;
    input [4:0] input_805;
    input [4:0] input_806;
    input [4:0] input_807;
    input [4:0] input_808;
    input [4:0] input_809;
    input [4:0] input_810;
    input [4:0] input_811;
    input [4:0] input_812;
    input [4:0] input_813;
    input [4:0] input_814;
    input [4:0] input_815;
    input [4:0] input_816;
    input [4:0] input_817;
    input [4:0] input_818;
    input [4:0] input_819;
    input [4:0] input_820;
    input [4:0] input_821;
    input [4:0] input_822;
    input [4:0] input_823;
    input [4:0] input_824;
    input [4:0] input_825;
    input [4:0] input_826;
    input [4:0] input_827;
    input [4:0] input_828;
    input [4:0] input_829;
    input [4:0] input_830;
    input [4:0] input_831;
    input [4:0] input_832;
    input [4:0] input_833;
    input [4:0] input_834;
    input [4:0] input_835;
    input [4:0] input_836;
    input [4:0] input_837;
    input [4:0] input_838;
    input [4:0] input_839;
    input [4:0] input_840;
    input [4:0] input_841;
    input [4:0] input_842;
    input [4:0] input_843;
    input [4:0] input_844;
    input [4:0] input_845;
    input [4:0] input_846;
    input [4:0] input_847;
    input [4:0] input_848;
    input [4:0] input_849;
    input [4:0] input_850;
    input [4:0] input_851;
    input [4:0] input_852;
    input [4:0] input_853;
    input [4:0] input_854;
    input [4:0] input_855;
    input [4:0] input_856;
    input [4:0] input_857;
    input [4:0] input_858;
    input [4:0] input_859;
    input [4:0] input_860;
    input [4:0] input_861;
    input [4:0] input_862;
    input [4:0] input_863;
    input [4:0] input_864;
    input [4:0] input_865;
    input [4:0] input_866;
    input [4:0] input_867;
    input [4:0] input_868;
    input [4:0] input_869;
    input [4:0] input_870;
    input [4:0] input_871;
    input [4:0] input_872;
    input [4:0] input_873;
    input [4:0] input_874;
    input [4:0] input_875;
    input [4:0] input_876;
    input [4:0] input_877;
    input [4:0] input_878;
    input [4:0] input_879;
    input [4:0] input_880;
    input [4:0] input_881;
    input [4:0] input_882;
    input [4:0] input_883;
    input [4:0] input_884;
    input [4:0] input_885;
    input [4:0] input_886;
    input [4:0] input_887;
    input [4:0] input_888;
    input [4:0] input_889;
    input [4:0] input_890;
    input [4:0] input_891;
    input [4:0] input_892;
    input [4:0] input_893;
    input [4:0] input_894;
    input [4:0] input_895;
    input [4:0] input_896;
    input [4:0] input_897;
    input [4:0] input_898;
    input [4:0] input_899;
    input [4:0] input_900;
    input [4:0] input_901;
    input [4:0] input_902;
    input [4:0] input_903;
    input [4:0] input_904;
    input [4:0] input_905;
    input [4:0] input_906;
    input [4:0] input_907;
    input [4:0] input_908;
    input [4:0] input_909;
    input [4:0] input_910;
    input [4:0] input_911;
    input [4:0] input_912;
    input [4:0] input_913;
    input [4:0] input_914;
    input [4:0] input_915;
    input [4:0] input_916;
    input [4:0] input_917;
    input [4:0] input_918;
    input [4:0] input_919;
    input [4:0] input_920;
    input [4:0] input_921;
    input [4:0] input_922;
    input [4:0] input_923;
    input [4:0] input_924;
    input [4:0] input_925;
    input [4:0] input_926;
    input [4:0] input_927;
    input [4:0] input_928;
    input [4:0] input_929;
    input [4:0] input_930;
    input [4:0] input_931;
    input [4:0] input_932;
    input [4:0] input_933;
    input [4:0] input_934;
    input [4:0] input_935;
    input [4:0] input_936;
    input [4:0] input_937;
    input [4:0] input_938;
    input [4:0] input_939;
    input [4:0] input_940;
    input [4:0] input_941;
    input [4:0] input_942;
    input [4:0] input_943;
    input [4:0] input_944;
    input [4:0] input_945;
    input [4:0] input_946;
    input [4:0] input_947;
    input [4:0] input_948;
    input [4:0] input_949;
    input [4:0] input_950;
    input [4:0] input_951;
    input [4:0] input_952;
    input [4:0] input_953;
    input [4:0] input_954;
    input [4:0] input_955;
    input [4:0] input_956;
    input [4:0] input_957;
    input [4:0] input_958;
    input [4:0] input_959;
    input [4:0] input_960;
    input [4:0] input_961;
    input [4:0] input_962;
    input [4:0] input_963;
    input [4:0] input_964;
    input [4:0] input_965;
    input [4:0] input_966;
    input [4:0] input_967;
    input [4:0] input_968;
    input [4:0] input_969;
    input [4:0] input_970;
    input [4:0] input_971;
    input [4:0] input_972;
    input [4:0] input_973;
    input [4:0] input_974;
    input [4:0] input_975;
    input [4:0] input_976;
    input [4:0] input_977;
    input [4:0] input_978;
    input [4:0] input_979;
    input [4:0] input_980;
    input [4:0] input_981;
    input [4:0] input_982;
    input [4:0] input_983;
    input [4:0] input_984;
    input [4:0] input_985;
    input [4:0] input_986;
    input [4:0] input_987;
    input [4:0] input_988;
    input [4:0] input_989;
    input [4:0] input_990;
    input [4:0] input_991;
    input [4:0] input_992;
    input [4:0] input_993;
    input [4:0] input_994;
    input [4:0] input_995;
    input [4:0] input_996;
    input [4:0] input_997;
    input [4:0] input_998;
    input [4:0] input_999;
    input [4:0] input_1000;
    input [4:0] input_1001;
    input [4:0] input_1002;
    input [4:0] input_1003;
    input [4:0] input_1004;
    input [4:0] input_1005;
    input [4:0] input_1006;
    input [4:0] input_1007;
    input [4:0] input_1008;
    input [4:0] input_1009;
    input [4:0] input_1010;
    input [4:0] input_1011;
    input [4:0] input_1012;
    input [4:0] input_1013;
    input [4:0] input_1014;
    input [4:0] input_1015;
    input [4:0] input_1016;
    input [4:0] input_1017;
    input [4:0] input_1018;
    input [4:0] input_1019;
    input [4:0] input_1020;
    input [4:0] input_1021;
    input [4:0] input_1022;
    input [4:0] input_1023;
    input [4:0] input_1024;
    input [4:0] input_1025;
    input [4:0] input_1026;
    input [4:0] input_1027;
    input [4:0] input_1028;
    input [4:0] input_1029;
    input [4:0] input_1030;
    input [4:0] input_1031;
    input [4:0] input_1032;
    input [4:0] input_1033;
    input [4:0] input_1034;
    input [4:0] input_1035;
    input [4:0] input_1036;
    input [4:0] input_1037;
    input [4:0] input_1038;
    input [4:0] input_1039;
    input [4:0] input_1040;
    input [4:0] input_1041;
    input [4:0] input_1042;
    input [4:0] input_1043;
    input [4:0] input_1044;
    input [4:0] input_1045;
    input [4:0] input_1046;
    input [4:0] input_1047;
    input [4:0] input_1048;
    input [4:0] input_1049;
    input [4:0] input_1050;
    input [4:0] input_1051;
    input [4:0] input_1052;
    input [4:0] input_1053;
    input [4:0] input_1054;
    input [4:0] input_1055;
    input [4:0] input_1056;
    input [4:0] input_1057;
    input [4:0] input_1058;
    input [4:0] input_1059;
    input [4:0] input_1060;
    input [4:0] input_1061;
    input [4:0] input_1062;
    input [4:0] input_1063;
    input [4:0] input_1064;
    input [4:0] input_1065;
    input [4:0] input_1066;
    input [4:0] input_1067;
    input [4:0] input_1068;
    input [4:0] input_1069;
    input [4:0] input_1070;
    input [4:0] input_1071;
    input [4:0] input_1072;
    input [4:0] input_1073;
    input [4:0] input_1074;
    input [4:0] input_1075;
    input [4:0] input_1076;
    input [4:0] input_1077;
    input [4:0] input_1078;
    input [4:0] input_1079;
    input [4:0] input_1080;
    input [4:0] input_1081;
    input [4:0] input_1082;
    input [4:0] input_1083;
    input [4:0] input_1084;
    input [4:0] input_1085;
    input [4:0] input_1086;
    input [4:0] input_1087;
    input [4:0] input_1088;
    input [4:0] input_1089;
    input [4:0] input_1090;
    input [4:0] input_1091;
    input [4:0] input_1092;
    input [4:0] input_1093;
    input [4:0] input_1094;
    input [4:0] input_1095;
    input [4:0] input_1096;
    input [4:0] input_1097;
    input [4:0] input_1098;
    input [4:0] input_1099;
    input [4:0] input_1100;
    input [4:0] input_1101;
    input [4:0] input_1102;
    input [4:0] input_1103;
    input [4:0] input_1104;
    input [4:0] input_1105;
    input [4:0] input_1106;
    input [4:0] input_1107;
    input [4:0] input_1108;
    input [4:0] input_1109;
    input [4:0] input_1110;
    input [4:0] input_1111;
    input [4:0] input_1112;
    input [4:0] input_1113;
    input [4:0] input_1114;
    input [4:0] input_1115;
    input [4:0] input_1116;
    input [4:0] input_1117;
    input [4:0] input_1118;
    input [4:0] input_1119;
    input [4:0] input_1120;
    input [4:0] input_1121;
    input [4:0] input_1122;
    input [4:0] input_1123;
    input [4:0] input_1124;
    input [4:0] input_1125;
    input [4:0] input_1126;
    input [4:0] input_1127;
    input [4:0] input_1128;
    input [4:0] input_1129;
    input [4:0] input_1130;
    input [4:0] input_1131;
    input [4:0] input_1132;
    input [4:0] input_1133;
    input [4:0] input_1134;
    input [4:0] input_1135;
    input [4:0] input_1136;
    input [4:0] input_1137;
    input [4:0] input_1138;
    input [4:0] input_1139;
    input [4:0] input_1140;
    input [4:0] input_1141;
    input [4:0] input_1142;
    input [4:0] input_1143;
    input [4:0] input_1144;
    input [4:0] input_1145;
    input [4:0] input_1146;
    input [4:0] input_1147;
    input [4:0] input_1148;
    input [4:0] input_1149;
    input [4:0] input_1150;
    input [4:0] input_1151;
    input [4:0] input_1152;
    input [4:0] input_1153;
    input [4:0] input_1154;
    input [4:0] input_1155;
    input [4:0] input_1156;
    input [4:0] input_1157;
    input [4:0] input_1158;
    input [4:0] input_1159;
    input [4:0] input_1160;
    input [4:0] input_1161;
    input [4:0] input_1162;
    input [4:0] input_1163;
    input [4:0] input_1164;
    input [4:0] input_1165;
    input [4:0] input_1166;
    input [4:0] input_1167;
    input [4:0] input_1168;
    input [4:0] input_1169;
    input [4:0] input_1170;
    input [4:0] input_1171;
    input [4:0] input_1172;
    input [4:0] input_1173;
    input [4:0] input_1174;
    input [4:0] input_1175;
    input [4:0] input_1176;
    input [4:0] input_1177;
    input [4:0] input_1178;
    input [4:0] input_1179;
    input [4:0] input_1180;
    input [4:0] input_1181;
    input [4:0] input_1182;
    input [4:0] input_1183;
    input [4:0] input_1184;
    input [4:0] input_1185;
    input [4:0] input_1186;
    input [4:0] input_1187;
    input [4:0] input_1188;
    input [4:0] input_1189;
    input [4:0] input_1190;
    input [4:0] input_1191;
    input [4:0] input_1192;
    input [4:0] input_1193;
    input [4:0] input_1194;
    input [4:0] input_1195;
    input [4:0] input_1196;
    input [4:0] input_1197;
    input [4:0] input_1198;
    input [4:0] input_1199;
    input [4:0] input_1200;
    input [4:0] input_1201;
    input [4:0] input_1202;
    input [4:0] input_1203;
    input [4:0] input_1204;
    input [4:0] input_1205;
    input [4:0] input_1206;
    input [4:0] input_1207;
    input [4:0] input_1208;
    input [4:0] input_1209;
    input [4:0] input_1210;
    input [4:0] input_1211;
    input [4:0] input_1212;
    input [4:0] input_1213;
    input [4:0] input_1214;
    input [4:0] input_1215;
    input [4:0] input_1216;
    input [4:0] input_1217;
    input [4:0] input_1218;
    input [4:0] input_1219;
    input [4:0] input_1220;
    input [4:0] input_1221;
    input [4:0] input_1222;
    input [4:0] input_1223;
    input [4:0] input_1224;
    input [4:0] input_1225;
    input [4:0] input_1226;
    input [4:0] input_1227;
    input [4:0] input_1228;
    input [4:0] input_1229;
    input [4:0] input_1230;
    input [4:0] input_1231;
    input [4:0] input_1232;
    input [4:0] input_1233;
    input [4:0] input_1234;
    input [4:0] input_1235;
    input [4:0] input_1236;
    input [4:0] input_1237;
    input [4:0] input_1238;
    input [4:0] input_1239;
    input [4:0] input_1240;
    input [4:0] input_1241;
    input [4:0] input_1242;
    input [4:0] input_1243;
    input [4:0] input_1244;
    input [4:0] input_1245;
    input [4:0] input_1246;
    input [4:0] input_1247;
    input [4:0] input_1248;
    input [4:0] input_1249;
    input [4:0] input_1250;
    input [4:0] input_1251;
    input [4:0] input_1252;
    input [4:0] input_1253;
    input [4:0] input_1254;
    input [4:0] input_1255;
    input [4:0] input_1256;
    input [4:0] input_1257;
    input [4:0] input_1258;
    input [4:0] input_1259;
    input [4:0] input_1260;
    input [4:0] input_1261;
    input [4:0] input_1262;
    input [4:0] input_1263;
    input [4:0] input_1264;
    input [4:0] input_1265;
    input [4:0] input_1266;
    input [4:0] input_1267;
    input [4:0] input_1268;
    input [4:0] input_1269;
    input [4:0] input_1270;
    input [4:0] input_1271;
    input [4:0] input_1272;
    input [4:0] input_1273;
    input [4:0] input_1274;
    input [4:0] input_1275;
    input [4:0] input_1276;
    input [4:0] input_1277;
    input [4:0] input_1278;
    input [4:0] input_1279;
    input [4:0] input_1280;
    input [4:0] input_1281;
    input [4:0] input_1282;
    input [4:0] input_1283;
    input [4:0] input_1284;
    input [4:0] input_1285;
    input [4:0] input_1286;
    input [4:0] input_1287;
    input [4:0] input_1288;
    input [4:0] input_1289;
    input [4:0] input_1290;
    input [4:0] input_1291;
    input [4:0] input_1292;
    input [4:0] input_1293;
    input [4:0] input_1294;
    input [4:0] input_1295;
    input [4:0] input_1296;
    input [4:0] input_1297;
    input [4:0] input_1298;
    input [4:0] input_1299;
    input [4:0] input_1300;
    input [4:0] input_1301;
    input [4:0] input_1302;
    input [4:0] input_1303;
    input [4:0] input_1304;
    input [4:0] input_1305;
    input [4:0] input_1306;
    input [4:0] input_1307;
    input [4:0] input_1308;
    input [4:0] input_1309;
    input [4:0] input_1310;
    input [4:0] input_1311;
    input [4:0] input_1312;
    input [4:0] input_1313;
    input [4:0] input_1314;
    input [4:0] input_1315;
    input [4:0] input_1316;
    input [4:0] input_1317;
    input [4:0] input_1318;
    input [4:0] input_1319;
    input [4:0] input_1320;
    input [4:0] input_1321;
    input [4:0] input_1322;
    input [4:0] input_1323;
    input [4:0] input_1324;
    input [4:0] input_1325;
    input [4:0] input_1326;
    input [4:0] input_1327;
    input [4:0] input_1328;
    input [4:0] input_1329;
    input [4:0] input_1330;
    input [4:0] input_1331;
    input [4:0] input_1332;
    input [4:0] input_1333;
    input [4:0] input_1334;
    input [4:0] input_1335;
    input [4:0] input_1336;
    input [4:0] input_1337;
    input [4:0] input_1338;
    input [4:0] input_1339;
    input [4:0] input_1340;
    input [4:0] input_1341;
    input [4:0] input_1342;
    input [4:0] input_1343;
    input [4:0] input_1344;
    input [4:0] input_1345;
    input [4:0] input_1346;
    input [4:0] input_1347;
    input [4:0] input_1348;
    input [4:0] input_1349;
    input [4:0] input_1350;
    input [4:0] input_1351;
    input [4:0] input_1352;
    input [4:0] input_1353;
    input [4:0] input_1354;
    input [4:0] input_1355;
    input [4:0] input_1356;
    input [4:0] input_1357;
    input [4:0] input_1358;
    input [4:0] input_1359;
    input [4:0] input_1360;
    input [4:0] input_1361;
    input [4:0] input_1362;
    input [4:0] input_1363;
    input [4:0] input_1364;
    input [4:0] input_1365;
    input [4:0] input_1366;
    input [4:0] input_1367;
    input [4:0] input_1368;
    input [4:0] input_1369;
    input [4:0] input_1370;
    input [4:0] input_1371;
    input [4:0] input_1372;
    input [4:0] input_1373;
    input [4:0] input_1374;
    input [4:0] input_1375;
    input [4:0] input_1376;
    input [4:0] input_1377;
    input [4:0] input_1378;
    input [4:0] input_1379;
    input [4:0] input_1380;
    input [4:0] input_1381;
    input [4:0] input_1382;
    input [4:0] input_1383;
    input [4:0] input_1384;
    input [4:0] input_1385;
    input [4:0] input_1386;
    input [4:0] input_1387;
    input [4:0] input_1388;
    input [4:0] input_1389;
    input [4:0] input_1390;
    input [4:0] input_1391;
    input [4:0] input_1392;
    input [4:0] input_1393;
    input [4:0] input_1394;
    input [4:0] input_1395;
    input [4:0] input_1396;
    input [4:0] input_1397;
    input [4:0] input_1398;
    input [4:0] input_1399;
    input [4:0] input_1400;
    input [4:0] input_1401;
    input [4:0] input_1402;
    input [4:0] input_1403;
    input [4:0] input_1404;
    input [4:0] input_1405;
    input [4:0] input_1406;
    input [4:0] input_1407;
    input [4:0] input_1408;
    input [4:0] input_1409;
    input [4:0] input_1410;
    input [4:0] input_1411;
    input [4:0] input_1412;
    input [4:0] input_1413;
    input [4:0] input_1414;
    input [4:0] input_1415;
    input [4:0] input_1416;
    input [4:0] input_1417;
    input [4:0] input_1418;
    input [4:0] input_1419;
    input [4:0] input_1420;
    input [4:0] input_1421;
    input [4:0] input_1422;
    input [4:0] input_1423;
    input [4:0] input_1424;
    input [4:0] input_1425;
    input [4:0] input_1426;
    input [4:0] input_1427;
    input [4:0] input_1428;
    input [4:0] input_1429;
    input [4:0] input_1430;
    input [4:0] input_1431;
    input [4:0] input_1432;
    input [4:0] input_1433;
    input [4:0] input_1434;
    input [4:0] input_1435;
    input [4:0] input_1436;
    input [4:0] input_1437;
    input [4:0] input_1438;
    input [4:0] input_1439;
    input [4:0] input_1440;
    input [4:0] input_1441;
    input [4:0] input_1442;
    input [4:0] input_1443;
    input [4:0] input_1444;
    input [4:0] input_1445;
    input [4:0] input_1446;
    input [4:0] input_1447;
    input [4:0] input_1448;
    input [4:0] input_1449;
    input [4:0] input_1450;
    input [4:0] input_1451;
    input [4:0] input_1452;
    input [4:0] input_1453;
    input [4:0] input_1454;
    input [4:0] input_1455;
    input [4:0] input_1456;
    input [4:0] input_1457;
    input [4:0] input_1458;
    input [4:0] input_1459;
    input [4:0] input_1460;
    input [4:0] input_1461;
    input [4:0] input_1462;
    input [4:0] input_1463;
    input [4:0] input_1464;
    input [4:0] input_1465;
    input [4:0] input_1466;
    input [4:0] input_1467;
    input [4:0] input_1468;
    input [4:0] input_1469;
    input [4:0] input_1470;
    input [4:0] input_1471;
    input [4:0] input_1472;
    input [4:0] input_1473;
    input [4:0] input_1474;
    input [4:0] input_1475;
    input [4:0] input_1476;
    input [4:0] input_1477;
    input [4:0] input_1478;
    input [4:0] input_1479;
    input [4:0] input_1480;
    input [4:0] input_1481;
    input [4:0] input_1482;
    input [4:0] input_1483;
    input [4:0] input_1484;
    input [4:0] input_1485;
    input [4:0] input_1486;
    input [4:0] input_1487;
    input [4:0] input_1488;
    input [4:0] input_1489;
    input [4:0] input_1490;
    input [4:0] input_1491;
    input [4:0] input_1492;
    input [4:0] input_1493;
    input [4:0] input_1494;
    input [4:0] input_1495;
    input [4:0] input_1496;
    input [4:0] input_1497;
    input [4:0] input_1498;
    input [4:0] input_1499;
    input [4:0] input_1500;
    input [4:0] input_1501;
    input [4:0] input_1502;
    input [4:0] input_1503;
    input [4:0] input_1504;
    input [4:0] input_1505;
    input [4:0] input_1506;
    input [4:0] input_1507;
    input [4:0] input_1508;
    input [4:0] input_1509;
    input [4:0] input_1510;
    input [4:0] input_1511;
    input [4:0] input_1512;
    input [4:0] input_1513;
    input [4:0] input_1514;
    input [4:0] input_1515;
    input [4:0] input_1516;
    input [4:0] input_1517;
    input [4:0] input_1518;
    input [4:0] input_1519;
    input [4:0] input_1520;
    input [4:0] input_1521;
    input [4:0] input_1522;
    input [4:0] input_1523;
    input [4:0] input_1524;
    input [4:0] input_1525;
    input [4:0] input_1526;
    input [4:0] input_1527;
    input [4:0] input_1528;
    input [4:0] input_1529;
    input [4:0] input_1530;
    input [4:0] input_1531;
    input [4:0] input_1532;
    input [4:0] input_1533;
    input [4:0] input_1534;
    input [4:0] input_1535;
    input [4:0] input_1536;
    input [4:0] input_1537;
    input [4:0] input_1538;
    input [4:0] input_1539;
    input [4:0] input_1540;
    input [4:0] input_1541;
    input [4:0] input_1542;
    input [4:0] input_1543;
    input [4:0] input_1544;
    input [4:0] input_1545;
    input [4:0] input_1546;
    input [4:0] input_1547;
    input [4:0] input_1548;
    input [4:0] input_1549;
    input [4:0] input_1550;
    input [4:0] input_1551;
    input [4:0] input_1552;
    input [4:0] input_1553;
    input [4:0] input_1554;
    input [4:0] input_1555;
    input [4:0] input_1556;
    input [4:0] input_1557;
    input [4:0] input_1558;
    input [4:0] input_1559;
    input [4:0] input_1560;
    input [4:0] input_1561;
    input [4:0] input_1562;
    input [4:0] input_1563;
    input [4:0] input_1564;
    input [4:0] input_1565;
    input [4:0] input_1566;
    input [4:0] input_1567;
    input [4:0] input_1568;
    input [4:0] input_1569;
    input [4:0] input_1570;
    input [4:0] input_1571;
    input [4:0] input_1572;
    input [4:0] input_1573;
    input [4:0] input_1574;
    input [4:0] input_1575;
    input [4:0] input_1576;
    input [4:0] input_1577;
    input [4:0] input_1578;
    input [4:0] input_1579;
    input [4:0] input_1580;
    input [4:0] input_1581;
    input [4:0] input_1582;
    input [4:0] input_1583;
    input [4:0] input_1584;
    input [4:0] input_1585;
    input [4:0] input_1586;
    input [4:0] input_1587;
    input [4:0] input_1588;
    input [4:0] input_1589;
    input [4:0] input_1590;
    input [4:0] input_1591;
    input [4:0] input_1592;
    input [4:0] input_1593;
    input [4:0] input_1594;
    input [4:0] input_1595;
    input [4:0] input_1596;
    input [4:0] input_1597;
    input [4:0] input_1598;
    input [4:0] input_1599;
    input [4:0] input_1600;
    input [4:0] input_1601;
    input [4:0] input_1602;
    input [4:0] input_1603;
    input [4:0] input_1604;
    input [4:0] input_1605;
    input [4:0] input_1606;
    input [4:0] input_1607;
    input [4:0] input_1608;
    input [4:0] input_1609;
    input [4:0] input_1610;
    input [4:0] input_1611;
    input [4:0] input_1612;
    input [4:0] input_1613;
    input [4:0] input_1614;
    input [4:0] input_1615;
    input [4:0] input_1616;
    input [4:0] input_1617;
    input [4:0] input_1618;
    input [4:0] input_1619;
    input [4:0] input_1620;
    input [4:0] input_1621;
    input [4:0] input_1622;
    input [4:0] input_1623;
    input [4:0] input_1624;
    input [4:0] input_1625;
    input [4:0] input_1626;
    input [4:0] input_1627;
    input [4:0] input_1628;
    input [4:0] input_1629;
    input [4:0] input_1630;
    input [4:0] input_1631;
    input [4:0] input_1632;
    input [4:0] input_1633;
    input [4:0] input_1634;
    input [4:0] input_1635;
    input [4:0] input_1636;
    input [4:0] input_1637;
    input [4:0] input_1638;
    input [4:0] input_1639;
    input [4:0] input_1640;
    input [4:0] input_1641;
    input [4:0] input_1642;
    input [4:0] input_1643;
    input [4:0] input_1644;
    input [4:0] input_1645;
    input [4:0] input_1646;
    input [4:0] input_1647;
    input [4:0] input_1648;
    input [4:0] input_1649;
    input [4:0] input_1650;
    input [4:0] input_1651;
    input [4:0] input_1652;
    input [4:0] input_1653;
    input [4:0] input_1654;
    input [4:0] input_1655;
    input [4:0] input_1656;
    input [4:0] input_1657;
    input [4:0] input_1658;
    input [4:0] input_1659;
    input [4:0] input_1660;
    input [4:0] input_1661;
    input [4:0] input_1662;
    input [4:0] input_1663;
    input [4:0] input_1664;
    input [4:0] input_1665;
    input [4:0] input_1666;
    input [4:0] input_1667;
    input [4:0] input_1668;
    input [4:0] input_1669;
    input [4:0] input_1670;
    input [4:0] input_1671;
    input [4:0] input_1672;
    input [4:0] input_1673;
    input [4:0] input_1674;
    input [4:0] input_1675;
    input [4:0] input_1676;
    input [4:0] input_1677;
    input [4:0] input_1678;
    input [4:0] input_1679;
    input [4:0] input_1680;
    input [4:0] input_1681;
    input [4:0] input_1682;
    input [4:0] input_1683;
    input [4:0] input_1684;
    input [4:0] input_1685;
    input [4:0] input_1686;
    input [4:0] input_1687;
    input [4:0] input_1688;
    input [4:0] input_1689;
    input [4:0] input_1690;
    input [4:0] input_1691;
    input [4:0] input_1692;
    input [4:0] input_1693;
    input [4:0] input_1694;
    input [4:0] input_1695;
    input [4:0] input_1696;
    input [4:0] input_1697;
    input [4:0] input_1698;
    input [4:0] input_1699;
    input [4:0] input_1700;
    input [4:0] input_1701;
    input [4:0] input_1702;
    input [4:0] input_1703;
    input [4:0] input_1704;
    input [4:0] input_1705;
    input [4:0] input_1706;
    input [4:0] input_1707;
    input [4:0] input_1708;
    input [4:0] input_1709;
    input [4:0] input_1710;
    input [4:0] input_1711;
    input [4:0] input_1712;
    input [4:0] input_1713;
    input [4:0] input_1714;
    input [4:0] input_1715;
    input [4:0] input_1716;
    input [4:0] input_1717;
    input [4:0] input_1718;
    input [4:0] input_1719;
    input [4:0] input_1720;
    input [4:0] input_1721;
    input [4:0] input_1722;
    input [4:0] input_1723;
    input [4:0] input_1724;
    input [4:0] input_1725;
    input [4:0] input_1726;
    input [4:0] input_1727;
    input [4:0] input_1728;
    input [4:0] input_1729;
    input [4:0] input_1730;
    input [4:0] input_1731;
    input [4:0] input_1732;
    input [4:0] input_1733;
    input [4:0] input_1734;
    input [4:0] input_1735;
    input [4:0] input_1736;
    input [4:0] input_1737;
    input [4:0] input_1738;
    input [4:0] input_1739;
    input [4:0] input_1740;
    input [4:0] input_1741;
    input [4:0] input_1742;
    input [4:0] input_1743;
    input [4:0] input_1744;
    input [4:0] input_1745;
    input [4:0] input_1746;
    input [4:0] input_1747;
    input [4:0] input_1748;
    input [4:0] input_1749;
    input [4:0] input_1750;
    input [4:0] input_1751;
    input [4:0] input_1752;
    input [4:0] input_1753;
    input [4:0] input_1754;
    input [4:0] input_1755;
    input [4:0] input_1756;
    input [4:0] input_1757;
    input [4:0] input_1758;
    input [4:0] input_1759;
    input [4:0] input_1760;
    input [4:0] input_1761;
    input [4:0] input_1762;
    input [4:0] input_1763;
    input [4:0] input_1764;
    input [4:0] input_1765;
    input [4:0] input_1766;
    input [4:0] input_1767;
    input [4:0] input_1768;
    input [4:0] input_1769;
    input [4:0] input_1770;
    input [4:0] input_1771;
    input [4:0] input_1772;
    input [4:0] input_1773;
    input [4:0] input_1774;
    input [4:0] input_1775;
    input [4:0] input_1776;
    input [4:0] input_1777;
    input [4:0] input_1778;
    input [4:0] input_1779;
    input [4:0] input_1780;
    input [4:0] input_1781;
    input [4:0] input_1782;
    input [4:0] input_1783;
    input [4:0] input_1784;
    input [4:0] input_1785;
    input [4:0] input_1786;
    input [4:0] input_1787;
    input [4:0] input_1788;
    input [4:0] input_1789;
    input [4:0] input_1790;
    input [4:0] input_1791;
    input [10:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      11'b00000000000 : begin
        result = input_0;
      end
      11'b00000000001 : begin
        result = input_1;
      end
      11'b00000000010 : begin
        result = input_2;
      end
      11'b00000000011 : begin
        result = input_3;
      end
      11'b00000000100 : begin
        result = input_4;
      end
      11'b00000000101 : begin
        result = input_5;
      end
      11'b00000000110 : begin
        result = input_6;
      end
      11'b00000000111 : begin
        result = input_7;
      end
      11'b00000001000 : begin
        result = input_8;
      end
      11'b00000001001 : begin
        result = input_9;
      end
      11'b00000001010 : begin
        result = input_10;
      end
      11'b00000001011 : begin
        result = input_11;
      end
      11'b00000001100 : begin
        result = input_12;
      end
      11'b00000001101 : begin
        result = input_13;
      end
      11'b00000001110 : begin
        result = input_14;
      end
      11'b00000001111 : begin
        result = input_15;
      end
      11'b00000010000 : begin
        result = input_16;
      end
      11'b00000010001 : begin
        result = input_17;
      end
      11'b00000010010 : begin
        result = input_18;
      end
      11'b00000010011 : begin
        result = input_19;
      end
      11'b00000010100 : begin
        result = input_20;
      end
      11'b00000010101 : begin
        result = input_21;
      end
      11'b00000010110 : begin
        result = input_22;
      end
      11'b00000010111 : begin
        result = input_23;
      end
      11'b00000011000 : begin
        result = input_24;
      end
      11'b00000011001 : begin
        result = input_25;
      end
      11'b00000011010 : begin
        result = input_26;
      end
      11'b00000011011 : begin
        result = input_27;
      end
      11'b00000011100 : begin
        result = input_28;
      end
      11'b00000011101 : begin
        result = input_29;
      end
      11'b00000011110 : begin
        result = input_30;
      end
      11'b00000011111 : begin
        result = input_31;
      end
      11'b00000100000 : begin
        result = input_32;
      end
      11'b00000100001 : begin
        result = input_33;
      end
      11'b00000100010 : begin
        result = input_34;
      end
      11'b00000100011 : begin
        result = input_35;
      end
      11'b00000100100 : begin
        result = input_36;
      end
      11'b00000100101 : begin
        result = input_37;
      end
      11'b00000100110 : begin
        result = input_38;
      end
      11'b00000100111 : begin
        result = input_39;
      end
      11'b00000101000 : begin
        result = input_40;
      end
      11'b00000101001 : begin
        result = input_41;
      end
      11'b00000101010 : begin
        result = input_42;
      end
      11'b00000101011 : begin
        result = input_43;
      end
      11'b00000101100 : begin
        result = input_44;
      end
      11'b00000101101 : begin
        result = input_45;
      end
      11'b00000101110 : begin
        result = input_46;
      end
      11'b00000101111 : begin
        result = input_47;
      end
      11'b00000110000 : begin
        result = input_48;
      end
      11'b00000110001 : begin
        result = input_49;
      end
      11'b00000110010 : begin
        result = input_50;
      end
      11'b00000110011 : begin
        result = input_51;
      end
      11'b00000110100 : begin
        result = input_52;
      end
      11'b00000110101 : begin
        result = input_53;
      end
      11'b00000110110 : begin
        result = input_54;
      end
      11'b00000110111 : begin
        result = input_55;
      end
      11'b00000111000 : begin
        result = input_56;
      end
      11'b00000111001 : begin
        result = input_57;
      end
      11'b00000111010 : begin
        result = input_58;
      end
      11'b00000111011 : begin
        result = input_59;
      end
      11'b00000111100 : begin
        result = input_60;
      end
      11'b00000111101 : begin
        result = input_61;
      end
      11'b00000111110 : begin
        result = input_62;
      end
      11'b00000111111 : begin
        result = input_63;
      end
      11'b00001000000 : begin
        result = input_64;
      end
      11'b00001000001 : begin
        result = input_65;
      end
      11'b00001000010 : begin
        result = input_66;
      end
      11'b00001000011 : begin
        result = input_67;
      end
      11'b00001000100 : begin
        result = input_68;
      end
      11'b00001000101 : begin
        result = input_69;
      end
      11'b00001000110 : begin
        result = input_70;
      end
      11'b00001000111 : begin
        result = input_71;
      end
      11'b00001001000 : begin
        result = input_72;
      end
      11'b00001001001 : begin
        result = input_73;
      end
      11'b00001001010 : begin
        result = input_74;
      end
      11'b00001001011 : begin
        result = input_75;
      end
      11'b00001001100 : begin
        result = input_76;
      end
      11'b00001001101 : begin
        result = input_77;
      end
      11'b00001001110 : begin
        result = input_78;
      end
      11'b00001001111 : begin
        result = input_79;
      end
      11'b00001010000 : begin
        result = input_80;
      end
      11'b00001010001 : begin
        result = input_81;
      end
      11'b00001010010 : begin
        result = input_82;
      end
      11'b00001010011 : begin
        result = input_83;
      end
      11'b00001010100 : begin
        result = input_84;
      end
      11'b00001010101 : begin
        result = input_85;
      end
      11'b00001010110 : begin
        result = input_86;
      end
      11'b00001010111 : begin
        result = input_87;
      end
      11'b00001011000 : begin
        result = input_88;
      end
      11'b00001011001 : begin
        result = input_89;
      end
      11'b00001011010 : begin
        result = input_90;
      end
      11'b00001011011 : begin
        result = input_91;
      end
      11'b00001011100 : begin
        result = input_92;
      end
      11'b00001011101 : begin
        result = input_93;
      end
      11'b00001011110 : begin
        result = input_94;
      end
      11'b00001011111 : begin
        result = input_95;
      end
      11'b00001100000 : begin
        result = input_96;
      end
      11'b00001100001 : begin
        result = input_97;
      end
      11'b00001100010 : begin
        result = input_98;
      end
      11'b00001100011 : begin
        result = input_99;
      end
      11'b00001100100 : begin
        result = input_100;
      end
      11'b00001100101 : begin
        result = input_101;
      end
      11'b00001100110 : begin
        result = input_102;
      end
      11'b00001100111 : begin
        result = input_103;
      end
      11'b00001101000 : begin
        result = input_104;
      end
      11'b00001101001 : begin
        result = input_105;
      end
      11'b00001101010 : begin
        result = input_106;
      end
      11'b00001101011 : begin
        result = input_107;
      end
      11'b00001101100 : begin
        result = input_108;
      end
      11'b00001101101 : begin
        result = input_109;
      end
      11'b00001101110 : begin
        result = input_110;
      end
      11'b00001101111 : begin
        result = input_111;
      end
      11'b00001110000 : begin
        result = input_112;
      end
      11'b00001110001 : begin
        result = input_113;
      end
      11'b00001110010 : begin
        result = input_114;
      end
      11'b00001110011 : begin
        result = input_115;
      end
      11'b00001110100 : begin
        result = input_116;
      end
      11'b00001110101 : begin
        result = input_117;
      end
      11'b00001110110 : begin
        result = input_118;
      end
      11'b00001110111 : begin
        result = input_119;
      end
      11'b00001111000 : begin
        result = input_120;
      end
      11'b00001111001 : begin
        result = input_121;
      end
      11'b00001111010 : begin
        result = input_122;
      end
      11'b00001111011 : begin
        result = input_123;
      end
      11'b00001111100 : begin
        result = input_124;
      end
      11'b00001111101 : begin
        result = input_125;
      end
      11'b00001111110 : begin
        result = input_126;
      end
      11'b00001111111 : begin
        result = input_127;
      end
      11'b00010000000 : begin
        result = input_128;
      end
      11'b00010000001 : begin
        result = input_129;
      end
      11'b00010000010 : begin
        result = input_130;
      end
      11'b00010000011 : begin
        result = input_131;
      end
      11'b00010000100 : begin
        result = input_132;
      end
      11'b00010000101 : begin
        result = input_133;
      end
      11'b00010000110 : begin
        result = input_134;
      end
      11'b00010000111 : begin
        result = input_135;
      end
      11'b00010001000 : begin
        result = input_136;
      end
      11'b00010001001 : begin
        result = input_137;
      end
      11'b00010001010 : begin
        result = input_138;
      end
      11'b00010001011 : begin
        result = input_139;
      end
      11'b00010001100 : begin
        result = input_140;
      end
      11'b00010001101 : begin
        result = input_141;
      end
      11'b00010001110 : begin
        result = input_142;
      end
      11'b00010001111 : begin
        result = input_143;
      end
      11'b00010010000 : begin
        result = input_144;
      end
      11'b00010010001 : begin
        result = input_145;
      end
      11'b00010010010 : begin
        result = input_146;
      end
      11'b00010010011 : begin
        result = input_147;
      end
      11'b00010010100 : begin
        result = input_148;
      end
      11'b00010010101 : begin
        result = input_149;
      end
      11'b00010010110 : begin
        result = input_150;
      end
      11'b00010010111 : begin
        result = input_151;
      end
      11'b00010011000 : begin
        result = input_152;
      end
      11'b00010011001 : begin
        result = input_153;
      end
      11'b00010011010 : begin
        result = input_154;
      end
      11'b00010011011 : begin
        result = input_155;
      end
      11'b00010011100 : begin
        result = input_156;
      end
      11'b00010011101 : begin
        result = input_157;
      end
      11'b00010011110 : begin
        result = input_158;
      end
      11'b00010011111 : begin
        result = input_159;
      end
      11'b00010100000 : begin
        result = input_160;
      end
      11'b00010100001 : begin
        result = input_161;
      end
      11'b00010100010 : begin
        result = input_162;
      end
      11'b00010100011 : begin
        result = input_163;
      end
      11'b00010100100 : begin
        result = input_164;
      end
      11'b00010100101 : begin
        result = input_165;
      end
      11'b00010100110 : begin
        result = input_166;
      end
      11'b00010100111 : begin
        result = input_167;
      end
      11'b00010101000 : begin
        result = input_168;
      end
      11'b00010101001 : begin
        result = input_169;
      end
      11'b00010101010 : begin
        result = input_170;
      end
      11'b00010101011 : begin
        result = input_171;
      end
      11'b00010101100 : begin
        result = input_172;
      end
      11'b00010101101 : begin
        result = input_173;
      end
      11'b00010101110 : begin
        result = input_174;
      end
      11'b00010101111 : begin
        result = input_175;
      end
      11'b00010110000 : begin
        result = input_176;
      end
      11'b00010110001 : begin
        result = input_177;
      end
      11'b00010110010 : begin
        result = input_178;
      end
      11'b00010110011 : begin
        result = input_179;
      end
      11'b00010110100 : begin
        result = input_180;
      end
      11'b00010110101 : begin
        result = input_181;
      end
      11'b00010110110 : begin
        result = input_182;
      end
      11'b00010110111 : begin
        result = input_183;
      end
      11'b00010111000 : begin
        result = input_184;
      end
      11'b00010111001 : begin
        result = input_185;
      end
      11'b00010111010 : begin
        result = input_186;
      end
      11'b00010111011 : begin
        result = input_187;
      end
      11'b00010111100 : begin
        result = input_188;
      end
      11'b00010111101 : begin
        result = input_189;
      end
      11'b00010111110 : begin
        result = input_190;
      end
      11'b00010111111 : begin
        result = input_191;
      end
      11'b00011000000 : begin
        result = input_192;
      end
      11'b00011000001 : begin
        result = input_193;
      end
      11'b00011000010 : begin
        result = input_194;
      end
      11'b00011000011 : begin
        result = input_195;
      end
      11'b00011000100 : begin
        result = input_196;
      end
      11'b00011000101 : begin
        result = input_197;
      end
      11'b00011000110 : begin
        result = input_198;
      end
      11'b00011000111 : begin
        result = input_199;
      end
      11'b00011001000 : begin
        result = input_200;
      end
      11'b00011001001 : begin
        result = input_201;
      end
      11'b00011001010 : begin
        result = input_202;
      end
      11'b00011001011 : begin
        result = input_203;
      end
      11'b00011001100 : begin
        result = input_204;
      end
      11'b00011001101 : begin
        result = input_205;
      end
      11'b00011001110 : begin
        result = input_206;
      end
      11'b00011001111 : begin
        result = input_207;
      end
      11'b00011010000 : begin
        result = input_208;
      end
      11'b00011010001 : begin
        result = input_209;
      end
      11'b00011010010 : begin
        result = input_210;
      end
      11'b00011010011 : begin
        result = input_211;
      end
      11'b00011010100 : begin
        result = input_212;
      end
      11'b00011010101 : begin
        result = input_213;
      end
      11'b00011010110 : begin
        result = input_214;
      end
      11'b00011010111 : begin
        result = input_215;
      end
      11'b00011011000 : begin
        result = input_216;
      end
      11'b00011011001 : begin
        result = input_217;
      end
      11'b00011011010 : begin
        result = input_218;
      end
      11'b00011011011 : begin
        result = input_219;
      end
      11'b00011011100 : begin
        result = input_220;
      end
      11'b00011011101 : begin
        result = input_221;
      end
      11'b00011011110 : begin
        result = input_222;
      end
      11'b00011011111 : begin
        result = input_223;
      end
      11'b00011100000 : begin
        result = input_224;
      end
      11'b00011100001 : begin
        result = input_225;
      end
      11'b00011100010 : begin
        result = input_226;
      end
      11'b00011100011 : begin
        result = input_227;
      end
      11'b00011100100 : begin
        result = input_228;
      end
      11'b00011100101 : begin
        result = input_229;
      end
      11'b00011100110 : begin
        result = input_230;
      end
      11'b00011100111 : begin
        result = input_231;
      end
      11'b00011101000 : begin
        result = input_232;
      end
      11'b00011101001 : begin
        result = input_233;
      end
      11'b00011101010 : begin
        result = input_234;
      end
      11'b00011101011 : begin
        result = input_235;
      end
      11'b00011101100 : begin
        result = input_236;
      end
      11'b00011101101 : begin
        result = input_237;
      end
      11'b00011101110 : begin
        result = input_238;
      end
      11'b00011101111 : begin
        result = input_239;
      end
      11'b00011110000 : begin
        result = input_240;
      end
      11'b00011110001 : begin
        result = input_241;
      end
      11'b00011110010 : begin
        result = input_242;
      end
      11'b00011110011 : begin
        result = input_243;
      end
      11'b00011110100 : begin
        result = input_244;
      end
      11'b00011110101 : begin
        result = input_245;
      end
      11'b00011110110 : begin
        result = input_246;
      end
      11'b00011110111 : begin
        result = input_247;
      end
      11'b00011111000 : begin
        result = input_248;
      end
      11'b00011111001 : begin
        result = input_249;
      end
      11'b00011111010 : begin
        result = input_250;
      end
      11'b00011111011 : begin
        result = input_251;
      end
      11'b00011111100 : begin
        result = input_252;
      end
      11'b00011111101 : begin
        result = input_253;
      end
      11'b00011111110 : begin
        result = input_254;
      end
      11'b00011111111 : begin
        result = input_255;
      end
      11'b00100000000 : begin
        result = input_256;
      end
      11'b00100000001 : begin
        result = input_257;
      end
      11'b00100000010 : begin
        result = input_258;
      end
      11'b00100000011 : begin
        result = input_259;
      end
      11'b00100000100 : begin
        result = input_260;
      end
      11'b00100000101 : begin
        result = input_261;
      end
      11'b00100000110 : begin
        result = input_262;
      end
      11'b00100000111 : begin
        result = input_263;
      end
      11'b00100001000 : begin
        result = input_264;
      end
      11'b00100001001 : begin
        result = input_265;
      end
      11'b00100001010 : begin
        result = input_266;
      end
      11'b00100001011 : begin
        result = input_267;
      end
      11'b00100001100 : begin
        result = input_268;
      end
      11'b00100001101 : begin
        result = input_269;
      end
      11'b00100001110 : begin
        result = input_270;
      end
      11'b00100001111 : begin
        result = input_271;
      end
      11'b00100010000 : begin
        result = input_272;
      end
      11'b00100010001 : begin
        result = input_273;
      end
      11'b00100010010 : begin
        result = input_274;
      end
      11'b00100010011 : begin
        result = input_275;
      end
      11'b00100010100 : begin
        result = input_276;
      end
      11'b00100010101 : begin
        result = input_277;
      end
      11'b00100010110 : begin
        result = input_278;
      end
      11'b00100010111 : begin
        result = input_279;
      end
      11'b00100011000 : begin
        result = input_280;
      end
      11'b00100011001 : begin
        result = input_281;
      end
      11'b00100011010 : begin
        result = input_282;
      end
      11'b00100011011 : begin
        result = input_283;
      end
      11'b00100011100 : begin
        result = input_284;
      end
      11'b00100011101 : begin
        result = input_285;
      end
      11'b00100011110 : begin
        result = input_286;
      end
      11'b00100011111 : begin
        result = input_287;
      end
      11'b00100100000 : begin
        result = input_288;
      end
      11'b00100100001 : begin
        result = input_289;
      end
      11'b00100100010 : begin
        result = input_290;
      end
      11'b00100100011 : begin
        result = input_291;
      end
      11'b00100100100 : begin
        result = input_292;
      end
      11'b00100100101 : begin
        result = input_293;
      end
      11'b00100100110 : begin
        result = input_294;
      end
      11'b00100100111 : begin
        result = input_295;
      end
      11'b00100101000 : begin
        result = input_296;
      end
      11'b00100101001 : begin
        result = input_297;
      end
      11'b00100101010 : begin
        result = input_298;
      end
      11'b00100101011 : begin
        result = input_299;
      end
      11'b00100101100 : begin
        result = input_300;
      end
      11'b00100101101 : begin
        result = input_301;
      end
      11'b00100101110 : begin
        result = input_302;
      end
      11'b00100101111 : begin
        result = input_303;
      end
      11'b00100110000 : begin
        result = input_304;
      end
      11'b00100110001 : begin
        result = input_305;
      end
      11'b00100110010 : begin
        result = input_306;
      end
      11'b00100110011 : begin
        result = input_307;
      end
      11'b00100110100 : begin
        result = input_308;
      end
      11'b00100110101 : begin
        result = input_309;
      end
      11'b00100110110 : begin
        result = input_310;
      end
      11'b00100110111 : begin
        result = input_311;
      end
      11'b00100111000 : begin
        result = input_312;
      end
      11'b00100111001 : begin
        result = input_313;
      end
      11'b00100111010 : begin
        result = input_314;
      end
      11'b00100111011 : begin
        result = input_315;
      end
      11'b00100111100 : begin
        result = input_316;
      end
      11'b00100111101 : begin
        result = input_317;
      end
      11'b00100111110 : begin
        result = input_318;
      end
      11'b00100111111 : begin
        result = input_319;
      end
      11'b00101000000 : begin
        result = input_320;
      end
      11'b00101000001 : begin
        result = input_321;
      end
      11'b00101000010 : begin
        result = input_322;
      end
      11'b00101000011 : begin
        result = input_323;
      end
      11'b00101000100 : begin
        result = input_324;
      end
      11'b00101000101 : begin
        result = input_325;
      end
      11'b00101000110 : begin
        result = input_326;
      end
      11'b00101000111 : begin
        result = input_327;
      end
      11'b00101001000 : begin
        result = input_328;
      end
      11'b00101001001 : begin
        result = input_329;
      end
      11'b00101001010 : begin
        result = input_330;
      end
      11'b00101001011 : begin
        result = input_331;
      end
      11'b00101001100 : begin
        result = input_332;
      end
      11'b00101001101 : begin
        result = input_333;
      end
      11'b00101001110 : begin
        result = input_334;
      end
      11'b00101001111 : begin
        result = input_335;
      end
      11'b00101010000 : begin
        result = input_336;
      end
      11'b00101010001 : begin
        result = input_337;
      end
      11'b00101010010 : begin
        result = input_338;
      end
      11'b00101010011 : begin
        result = input_339;
      end
      11'b00101010100 : begin
        result = input_340;
      end
      11'b00101010101 : begin
        result = input_341;
      end
      11'b00101010110 : begin
        result = input_342;
      end
      11'b00101010111 : begin
        result = input_343;
      end
      11'b00101011000 : begin
        result = input_344;
      end
      11'b00101011001 : begin
        result = input_345;
      end
      11'b00101011010 : begin
        result = input_346;
      end
      11'b00101011011 : begin
        result = input_347;
      end
      11'b00101011100 : begin
        result = input_348;
      end
      11'b00101011101 : begin
        result = input_349;
      end
      11'b00101011110 : begin
        result = input_350;
      end
      11'b00101011111 : begin
        result = input_351;
      end
      11'b00101100000 : begin
        result = input_352;
      end
      11'b00101100001 : begin
        result = input_353;
      end
      11'b00101100010 : begin
        result = input_354;
      end
      11'b00101100011 : begin
        result = input_355;
      end
      11'b00101100100 : begin
        result = input_356;
      end
      11'b00101100101 : begin
        result = input_357;
      end
      11'b00101100110 : begin
        result = input_358;
      end
      11'b00101100111 : begin
        result = input_359;
      end
      11'b00101101000 : begin
        result = input_360;
      end
      11'b00101101001 : begin
        result = input_361;
      end
      11'b00101101010 : begin
        result = input_362;
      end
      11'b00101101011 : begin
        result = input_363;
      end
      11'b00101101100 : begin
        result = input_364;
      end
      11'b00101101101 : begin
        result = input_365;
      end
      11'b00101101110 : begin
        result = input_366;
      end
      11'b00101101111 : begin
        result = input_367;
      end
      11'b00101110000 : begin
        result = input_368;
      end
      11'b00101110001 : begin
        result = input_369;
      end
      11'b00101110010 : begin
        result = input_370;
      end
      11'b00101110011 : begin
        result = input_371;
      end
      11'b00101110100 : begin
        result = input_372;
      end
      11'b00101110101 : begin
        result = input_373;
      end
      11'b00101110110 : begin
        result = input_374;
      end
      11'b00101110111 : begin
        result = input_375;
      end
      11'b00101111000 : begin
        result = input_376;
      end
      11'b00101111001 : begin
        result = input_377;
      end
      11'b00101111010 : begin
        result = input_378;
      end
      11'b00101111011 : begin
        result = input_379;
      end
      11'b00101111100 : begin
        result = input_380;
      end
      11'b00101111101 : begin
        result = input_381;
      end
      11'b00101111110 : begin
        result = input_382;
      end
      11'b00101111111 : begin
        result = input_383;
      end
      11'b00110000000 : begin
        result = input_384;
      end
      11'b00110000001 : begin
        result = input_385;
      end
      11'b00110000010 : begin
        result = input_386;
      end
      11'b00110000011 : begin
        result = input_387;
      end
      11'b00110000100 : begin
        result = input_388;
      end
      11'b00110000101 : begin
        result = input_389;
      end
      11'b00110000110 : begin
        result = input_390;
      end
      11'b00110000111 : begin
        result = input_391;
      end
      11'b00110001000 : begin
        result = input_392;
      end
      11'b00110001001 : begin
        result = input_393;
      end
      11'b00110001010 : begin
        result = input_394;
      end
      11'b00110001011 : begin
        result = input_395;
      end
      11'b00110001100 : begin
        result = input_396;
      end
      11'b00110001101 : begin
        result = input_397;
      end
      11'b00110001110 : begin
        result = input_398;
      end
      11'b00110001111 : begin
        result = input_399;
      end
      11'b00110010000 : begin
        result = input_400;
      end
      11'b00110010001 : begin
        result = input_401;
      end
      11'b00110010010 : begin
        result = input_402;
      end
      11'b00110010011 : begin
        result = input_403;
      end
      11'b00110010100 : begin
        result = input_404;
      end
      11'b00110010101 : begin
        result = input_405;
      end
      11'b00110010110 : begin
        result = input_406;
      end
      11'b00110010111 : begin
        result = input_407;
      end
      11'b00110011000 : begin
        result = input_408;
      end
      11'b00110011001 : begin
        result = input_409;
      end
      11'b00110011010 : begin
        result = input_410;
      end
      11'b00110011011 : begin
        result = input_411;
      end
      11'b00110011100 : begin
        result = input_412;
      end
      11'b00110011101 : begin
        result = input_413;
      end
      11'b00110011110 : begin
        result = input_414;
      end
      11'b00110011111 : begin
        result = input_415;
      end
      11'b00110100000 : begin
        result = input_416;
      end
      11'b00110100001 : begin
        result = input_417;
      end
      11'b00110100010 : begin
        result = input_418;
      end
      11'b00110100011 : begin
        result = input_419;
      end
      11'b00110100100 : begin
        result = input_420;
      end
      11'b00110100101 : begin
        result = input_421;
      end
      11'b00110100110 : begin
        result = input_422;
      end
      11'b00110100111 : begin
        result = input_423;
      end
      11'b00110101000 : begin
        result = input_424;
      end
      11'b00110101001 : begin
        result = input_425;
      end
      11'b00110101010 : begin
        result = input_426;
      end
      11'b00110101011 : begin
        result = input_427;
      end
      11'b00110101100 : begin
        result = input_428;
      end
      11'b00110101101 : begin
        result = input_429;
      end
      11'b00110101110 : begin
        result = input_430;
      end
      11'b00110101111 : begin
        result = input_431;
      end
      11'b00110110000 : begin
        result = input_432;
      end
      11'b00110110001 : begin
        result = input_433;
      end
      11'b00110110010 : begin
        result = input_434;
      end
      11'b00110110011 : begin
        result = input_435;
      end
      11'b00110110100 : begin
        result = input_436;
      end
      11'b00110110101 : begin
        result = input_437;
      end
      11'b00110110110 : begin
        result = input_438;
      end
      11'b00110110111 : begin
        result = input_439;
      end
      11'b00110111000 : begin
        result = input_440;
      end
      11'b00110111001 : begin
        result = input_441;
      end
      11'b00110111010 : begin
        result = input_442;
      end
      11'b00110111011 : begin
        result = input_443;
      end
      11'b00110111100 : begin
        result = input_444;
      end
      11'b00110111101 : begin
        result = input_445;
      end
      11'b00110111110 : begin
        result = input_446;
      end
      11'b00110111111 : begin
        result = input_447;
      end
      11'b00111000000 : begin
        result = input_448;
      end
      11'b00111000001 : begin
        result = input_449;
      end
      11'b00111000010 : begin
        result = input_450;
      end
      11'b00111000011 : begin
        result = input_451;
      end
      11'b00111000100 : begin
        result = input_452;
      end
      11'b00111000101 : begin
        result = input_453;
      end
      11'b00111000110 : begin
        result = input_454;
      end
      11'b00111000111 : begin
        result = input_455;
      end
      11'b00111001000 : begin
        result = input_456;
      end
      11'b00111001001 : begin
        result = input_457;
      end
      11'b00111001010 : begin
        result = input_458;
      end
      11'b00111001011 : begin
        result = input_459;
      end
      11'b00111001100 : begin
        result = input_460;
      end
      11'b00111001101 : begin
        result = input_461;
      end
      11'b00111001110 : begin
        result = input_462;
      end
      11'b00111001111 : begin
        result = input_463;
      end
      11'b00111010000 : begin
        result = input_464;
      end
      11'b00111010001 : begin
        result = input_465;
      end
      11'b00111010010 : begin
        result = input_466;
      end
      11'b00111010011 : begin
        result = input_467;
      end
      11'b00111010100 : begin
        result = input_468;
      end
      11'b00111010101 : begin
        result = input_469;
      end
      11'b00111010110 : begin
        result = input_470;
      end
      11'b00111010111 : begin
        result = input_471;
      end
      11'b00111011000 : begin
        result = input_472;
      end
      11'b00111011001 : begin
        result = input_473;
      end
      11'b00111011010 : begin
        result = input_474;
      end
      11'b00111011011 : begin
        result = input_475;
      end
      11'b00111011100 : begin
        result = input_476;
      end
      11'b00111011101 : begin
        result = input_477;
      end
      11'b00111011110 : begin
        result = input_478;
      end
      11'b00111011111 : begin
        result = input_479;
      end
      11'b00111100000 : begin
        result = input_480;
      end
      11'b00111100001 : begin
        result = input_481;
      end
      11'b00111100010 : begin
        result = input_482;
      end
      11'b00111100011 : begin
        result = input_483;
      end
      11'b00111100100 : begin
        result = input_484;
      end
      11'b00111100101 : begin
        result = input_485;
      end
      11'b00111100110 : begin
        result = input_486;
      end
      11'b00111100111 : begin
        result = input_487;
      end
      11'b00111101000 : begin
        result = input_488;
      end
      11'b00111101001 : begin
        result = input_489;
      end
      11'b00111101010 : begin
        result = input_490;
      end
      11'b00111101011 : begin
        result = input_491;
      end
      11'b00111101100 : begin
        result = input_492;
      end
      11'b00111101101 : begin
        result = input_493;
      end
      11'b00111101110 : begin
        result = input_494;
      end
      11'b00111101111 : begin
        result = input_495;
      end
      11'b00111110000 : begin
        result = input_496;
      end
      11'b00111110001 : begin
        result = input_497;
      end
      11'b00111110010 : begin
        result = input_498;
      end
      11'b00111110011 : begin
        result = input_499;
      end
      11'b00111110100 : begin
        result = input_500;
      end
      11'b00111110101 : begin
        result = input_501;
      end
      11'b00111110110 : begin
        result = input_502;
      end
      11'b00111110111 : begin
        result = input_503;
      end
      11'b00111111000 : begin
        result = input_504;
      end
      11'b00111111001 : begin
        result = input_505;
      end
      11'b00111111010 : begin
        result = input_506;
      end
      11'b00111111011 : begin
        result = input_507;
      end
      11'b00111111100 : begin
        result = input_508;
      end
      11'b00111111101 : begin
        result = input_509;
      end
      11'b00111111110 : begin
        result = input_510;
      end
      11'b00111111111 : begin
        result = input_511;
      end
      11'b01000000000 : begin
        result = input_512;
      end
      11'b01000000001 : begin
        result = input_513;
      end
      11'b01000000010 : begin
        result = input_514;
      end
      11'b01000000011 : begin
        result = input_515;
      end
      11'b01000000100 : begin
        result = input_516;
      end
      11'b01000000101 : begin
        result = input_517;
      end
      11'b01000000110 : begin
        result = input_518;
      end
      11'b01000000111 : begin
        result = input_519;
      end
      11'b01000001000 : begin
        result = input_520;
      end
      11'b01000001001 : begin
        result = input_521;
      end
      11'b01000001010 : begin
        result = input_522;
      end
      11'b01000001011 : begin
        result = input_523;
      end
      11'b01000001100 : begin
        result = input_524;
      end
      11'b01000001101 : begin
        result = input_525;
      end
      11'b01000001110 : begin
        result = input_526;
      end
      11'b01000001111 : begin
        result = input_527;
      end
      11'b01000010000 : begin
        result = input_528;
      end
      11'b01000010001 : begin
        result = input_529;
      end
      11'b01000010010 : begin
        result = input_530;
      end
      11'b01000010011 : begin
        result = input_531;
      end
      11'b01000010100 : begin
        result = input_532;
      end
      11'b01000010101 : begin
        result = input_533;
      end
      11'b01000010110 : begin
        result = input_534;
      end
      11'b01000010111 : begin
        result = input_535;
      end
      11'b01000011000 : begin
        result = input_536;
      end
      11'b01000011001 : begin
        result = input_537;
      end
      11'b01000011010 : begin
        result = input_538;
      end
      11'b01000011011 : begin
        result = input_539;
      end
      11'b01000011100 : begin
        result = input_540;
      end
      11'b01000011101 : begin
        result = input_541;
      end
      11'b01000011110 : begin
        result = input_542;
      end
      11'b01000011111 : begin
        result = input_543;
      end
      11'b01000100000 : begin
        result = input_544;
      end
      11'b01000100001 : begin
        result = input_545;
      end
      11'b01000100010 : begin
        result = input_546;
      end
      11'b01000100011 : begin
        result = input_547;
      end
      11'b01000100100 : begin
        result = input_548;
      end
      11'b01000100101 : begin
        result = input_549;
      end
      11'b01000100110 : begin
        result = input_550;
      end
      11'b01000100111 : begin
        result = input_551;
      end
      11'b01000101000 : begin
        result = input_552;
      end
      11'b01000101001 : begin
        result = input_553;
      end
      11'b01000101010 : begin
        result = input_554;
      end
      11'b01000101011 : begin
        result = input_555;
      end
      11'b01000101100 : begin
        result = input_556;
      end
      11'b01000101101 : begin
        result = input_557;
      end
      11'b01000101110 : begin
        result = input_558;
      end
      11'b01000101111 : begin
        result = input_559;
      end
      11'b01000110000 : begin
        result = input_560;
      end
      11'b01000110001 : begin
        result = input_561;
      end
      11'b01000110010 : begin
        result = input_562;
      end
      11'b01000110011 : begin
        result = input_563;
      end
      11'b01000110100 : begin
        result = input_564;
      end
      11'b01000110101 : begin
        result = input_565;
      end
      11'b01000110110 : begin
        result = input_566;
      end
      11'b01000110111 : begin
        result = input_567;
      end
      11'b01000111000 : begin
        result = input_568;
      end
      11'b01000111001 : begin
        result = input_569;
      end
      11'b01000111010 : begin
        result = input_570;
      end
      11'b01000111011 : begin
        result = input_571;
      end
      11'b01000111100 : begin
        result = input_572;
      end
      11'b01000111101 : begin
        result = input_573;
      end
      11'b01000111110 : begin
        result = input_574;
      end
      11'b01000111111 : begin
        result = input_575;
      end
      11'b01001000000 : begin
        result = input_576;
      end
      11'b01001000001 : begin
        result = input_577;
      end
      11'b01001000010 : begin
        result = input_578;
      end
      11'b01001000011 : begin
        result = input_579;
      end
      11'b01001000100 : begin
        result = input_580;
      end
      11'b01001000101 : begin
        result = input_581;
      end
      11'b01001000110 : begin
        result = input_582;
      end
      11'b01001000111 : begin
        result = input_583;
      end
      11'b01001001000 : begin
        result = input_584;
      end
      11'b01001001001 : begin
        result = input_585;
      end
      11'b01001001010 : begin
        result = input_586;
      end
      11'b01001001011 : begin
        result = input_587;
      end
      11'b01001001100 : begin
        result = input_588;
      end
      11'b01001001101 : begin
        result = input_589;
      end
      11'b01001001110 : begin
        result = input_590;
      end
      11'b01001001111 : begin
        result = input_591;
      end
      11'b01001010000 : begin
        result = input_592;
      end
      11'b01001010001 : begin
        result = input_593;
      end
      11'b01001010010 : begin
        result = input_594;
      end
      11'b01001010011 : begin
        result = input_595;
      end
      11'b01001010100 : begin
        result = input_596;
      end
      11'b01001010101 : begin
        result = input_597;
      end
      11'b01001010110 : begin
        result = input_598;
      end
      11'b01001010111 : begin
        result = input_599;
      end
      11'b01001011000 : begin
        result = input_600;
      end
      11'b01001011001 : begin
        result = input_601;
      end
      11'b01001011010 : begin
        result = input_602;
      end
      11'b01001011011 : begin
        result = input_603;
      end
      11'b01001011100 : begin
        result = input_604;
      end
      11'b01001011101 : begin
        result = input_605;
      end
      11'b01001011110 : begin
        result = input_606;
      end
      11'b01001011111 : begin
        result = input_607;
      end
      11'b01001100000 : begin
        result = input_608;
      end
      11'b01001100001 : begin
        result = input_609;
      end
      11'b01001100010 : begin
        result = input_610;
      end
      11'b01001100011 : begin
        result = input_611;
      end
      11'b01001100100 : begin
        result = input_612;
      end
      11'b01001100101 : begin
        result = input_613;
      end
      11'b01001100110 : begin
        result = input_614;
      end
      11'b01001100111 : begin
        result = input_615;
      end
      11'b01001101000 : begin
        result = input_616;
      end
      11'b01001101001 : begin
        result = input_617;
      end
      11'b01001101010 : begin
        result = input_618;
      end
      11'b01001101011 : begin
        result = input_619;
      end
      11'b01001101100 : begin
        result = input_620;
      end
      11'b01001101101 : begin
        result = input_621;
      end
      11'b01001101110 : begin
        result = input_622;
      end
      11'b01001101111 : begin
        result = input_623;
      end
      11'b01001110000 : begin
        result = input_624;
      end
      11'b01001110001 : begin
        result = input_625;
      end
      11'b01001110010 : begin
        result = input_626;
      end
      11'b01001110011 : begin
        result = input_627;
      end
      11'b01001110100 : begin
        result = input_628;
      end
      11'b01001110101 : begin
        result = input_629;
      end
      11'b01001110110 : begin
        result = input_630;
      end
      11'b01001110111 : begin
        result = input_631;
      end
      11'b01001111000 : begin
        result = input_632;
      end
      11'b01001111001 : begin
        result = input_633;
      end
      11'b01001111010 : begin
        result = input_634;
      end
      11'b01001111011 : begin
        result = input_635;
      end
      11'b01001111100 : begin
        result = input_636;
      end
      11'b01001111101 : begin
        result = input_637;
      end
      11'b01001111110 : begin
        result = input_638;
      end
      11'b01001111111 : begin
        result = input_639;
      end
      11'b01010000000 : begin
        result = input_640;
      end
      11'b01010000001 : begin
        result = input_641;
      end
      11'b01010000010 : begin
        result = input_642;
      end
      11'b01010000011 : begin
        result = input_643;
      end
      11'b01010000100 : begin
        result = input_644;
      end
      11'b01010000101 : begin
        result = input_645;
      end
      11'b01010000110 : begin
        result = input_646;
      end
      11'b01010000111 : begin
        result = input_647;
      end
      11'b01010001000 : begin
        result = input_648;
      end
      11'b01010001001 : begin
        result = input_649;
      end
      11'b01010001010 : begin
        result = input_650;
      end
      11'b01010001011 : begin
        result = input_651;
      end
      11'b01010001100 : begin
        result = input_652;
      end
      11'b01010001101 : begin
        result = input_653;
      end
      11'b01010001110 : begin
        result = input_654;
      end
      11'b01010001111 : begin
        result = input_655;
      end
      11'b01010010000 : begin
        result = input_656;
      end
      11'b01010010001 : begin
        result = input_657;
      end
      11'b01010010010 : begin
        result = input_658;
      end
      11'b01010010011 : begin
        result = input_659;
      end
      11'b01010010100 : begin
        result = input_660;
      end
      11'b01010010101 : begin
        result = input_661;
      end
      11'b01010010110 : begin
        result = input_662;
      end
      11'b01010010111 : begin
        result = input_663;
      end
      11'b01010011000 : begin
        result = input_664;
      end
      11'b01010011001 : begin
        result = input_665;
      end
      11'b01010011010 : begin
        result = input_666;
      end
      11'b01010011011 : begin
        result = input_667;
      end
      11'b01010011100 : begin
        result = input_668;
      end
      11'b01010011101 : begin
        result = input_669;
      end
      11'b01010011110 : begin
        result = input_670;
      end
      11'b01010011111 : begin
        result = input_671;
      end
      11'b01010100000 : begin
        result = input_672;
      end
      11'b01010100001 : begin
        result = input_673;
      end
      11'b01010100010 : begin
        result = input_674;
      end
      11'b01010100011 : begin
        result = input_675;
      end
      11'b01010100100 : begin
        result = input_676;
      end
      11'b01010100101 : begin
        result = input_677;
      end
      11'b01010100110 : begin
        result = input_678;
      end
      11'b01010100111 : begin
        result = input_679;
      end
      11'b01010101000 : begin
        result = input_680;
      end
      11'b01010101001 : begin
        result = input_681;
      end
      11'b01010101010 : begin
        result = input_682;
      end
      11'b01010101011 : begin
        result = input_683;
      end
      11'b01010101100 : begin
        result = input_684;
      end
      11'b01010101101 : begin
        result = input_685;
      end
      11'b01010101110 : begin
        result = input_686;
      end
      11'b01010101111 : begin
        result = input_687;
      end
      11'b01010110000 : begin
        result = input_688;
      end
      11'b01010110001 : begin
        result = input_689;
      end
      11'b01010110010 : begin
        result = input_690;
      end
      11'b01010110011 : begin
        result = input_691;
      end
      11'b01010110100 : begin
        result = input_692;
      end
      11'b01010110101 : begin
        result = input_693;
      end
      11'b01010110110 : begin
        result = input_694;
      end
      11'b01010110111 : begin
        result = input_695;
      end
      11'b01010111000 : begin
        result = input_696;
      end
      11'b01010111001 : begin
        result = input_697;
      end
      11'b01010111010 : begin
        result = input_698;
      end
      11'b01010111011 : begin
        result = input_699;
      end
      11'b01010111100 : begin
        result = input_700;
      end
      11'b01010111101 : begin
        result = input_701;
      end
      11'b01010111110 : begin
        result = input_702;
      end
      11'b01010111111 : begin
        result = input_703;
      end
      11'b01011000000 : begin
        result = input_704;
      end
      11'b01011000001 : begin
        result = input_705;
      end
      11'b01011000010 : begin
        result = input_706;
      end
      11'b01011000011 : begin
        result = input_707;
      end
      11'b01011000100 : begin
        result = input_708;
      end
      11'b01011000101 : begin
        result = input_709;
      end
      11'b01011000110 : begin
        result = input_710;
      end
      11'b01011000111 : begin
        result = input_711;
      end
      11'b01011001000 : begin
        result = input_712;
      end
      11'b01011001001 : begin
        result = input_713;
      end
      11'b01011001010 : begin
        result = input_714;
      end
      11'b01011001011 : begin
        result = input_715;
      end
      11'b01011001100 : begin
        result = input_716;
      end
      11'b01011001101 : begin
        result = input_717;
      end
      11'b01011001110 : begin
        result = input_718;
      end
      11'b01011001111 : begin
        result = input_719;
      end
      11'b01011010000 : begin
        result = input_720;
      end
      11'b01011010001 : begin
        result = input_721;
      end
      11'b01011010010 : begin
        result = input_722;
      end
      11'b01011010011 : begin
        result = input_723;
      end
      11'b01011010100 : begin
        result = input_724;
      end
      11'b01011010101 : begin
        result = input_725;
      end
      11'b01011010110 : begin
        result = input_726;
      end
      11'b01011010111 : begin
        result = input_727;
      end
      11'b01011011000 : begin
        result = input_728;
      end
      11'b01011011001 : begin
        result = input_729;
      end
      11'b01011011010 : begin
        result = input_730;
      end
      11'b01011011011 : begin
        result = input_731;
      end
      11'b01011011100 : begin
        result = input_732;
      end
      11'b01011011101 : begin
        result = input_733;
      end
      11'b01011011110 : begin
        result = input_734;
      end
      11'b01011011111 : begin
        result = input_735;
      end
      11'b01011100000 : begin
        result = input_736;
      end
      11'b01011100001 : begin
        result = input_737;
      end
      11'b01011100010 : begin
        result = input_738;
      end
      11'b01011100011 : begin
        result = input_739;
      end
      11'b01011100100 : begin
        result = input_740;
      end
      11'b01011100101 : begin
        result = input_741;
      end
      11'b01011100110 : begin
        result = input_742;
      end
      11'b01011100111 : begin
        result = input_743;
      end
      11'b01011101000 : begin
        result = input_744;
      end
      11'b01011101001 : begin
        result = input_745;
      end
      11'b01011101010 : begin
        result = input_746;
      end
      11'b01011101011 : begin
        result = input_747;
      end
      11'b01011101100 : begin
        result = input_748;
      end
      11'b01011101101 : begin
        result = input_749;
      end
      11'b01011101110 : begin
        result = input_750;
      end
      11'b01011101111 : begin
        result = input_751;
      end
      11'b01011110000 : begin
        result = input_752;
      end
      11'b01011110001 : begin
        result = input_753;
      end
      11'b01011110010 : begin
        result = input_754;
      end
      11'b01011110011 : begin
        result = input_755;
      end
      11'b01011110100 : begin
        result = input_756;
      end
      11'b01011110101 : begin
        result = input_757;
      end
      11'b01011110110 : begin
        result = input_758;
      end
      11'b01011110111 : begin
        result = input_759;
      end
      11'b01011111000 : begin
        result = input_760;
      end
      11'b01011111001 : begin
        result = input_761;
      end
      11'b01011111010 : begin
        result = input_762;
      end
      11'b01011111011 : begin
        result = input_763;
      end
      11'b01011111100 : begin
        result = input_764;
      end
      11'b01011111101 : begin
        result = input_765;
      end
      11'b01011111110 : begin
        result = input_766;
      end
      11'b01011111111 : begin
        result = input_767;
      end
      11'b01100000000 : begin
        result = input_768;
      end
      11'b01100000001 : begin
        result = input_769;
      end
      11'b01100000010 : begin
        result = input_770;
      end
      11'b01100000011 : begin
        result = input_771;
      end
      11'b01100000100 : begin
        result = input_772;
      end
      11'b01100000101 : begin
        result = input_773;
      end
      11'b01100000110 : begin
        result = input_774;
      end
      11'b01100000111 : begin
        result = input_775;
      end
      11'b01100001000 : begin
        result = input_776;
      end
      11'b01100001001 : begin
        result = input_777;
      end
      11'b01100001010 : begin
        result = input_778;
      end
      11'b01100001011 : begin
        result = input_779;
      end
      11'b01100001100 : begin
        result = input_780;
      end
      11'b01100001101 : begin
        result = input_781;
      end
      11'b01100001110 : begin
        result = input_782;
      end
      11'b01100001111 : begin
        result = input_783;
      end
      11'b01100010000 : begin
        result = input_784;
      end
      11'b01100010001 : begin
        result = input_785;
      end
      11'b01100010010 : begin
        result = input_786;
      end
      11'b01100010011 : begin
        result = input_787;
      end
      11'b01100010100 : begin
        result = input_788;
      end
      11'b01100010101 : begin
        result = input_789;
      end
      11'b01100010110 : begin
        result = input_790;
      end
      11'b01100010111 : begin
        result = input_791;
      end
      11'b01100011000 : begin
        result = input_792;
      end
      11'b01100011001 : begin
        result = input_793;
      end
      11'b01100011010 : begin
        result = input_794;
      end
      11'b01100011011 : begin
        result = input_795;
      end
      11'b01100011100 : begin
        result = input_796;
      end
      11'b01100011101 : begin
        result = input_797;
      end
      11'b01100011110 : begin
        result = input_798;
      end
      11'b01100011111 : begin
        result = input_799;
      end
      11'b01100100000 : begin
        result = input_800;
      end
      11'b01100100001 : begin
        result = input_801;
      end
      11'b01100100010 : begin
        result = input_802;
      end
      11'b01100100011 : begin
        result = input_803;
      end
      11'b01100100100 : begin
        result = input_804;
      end
      11'b01100100101 : begin
        result = input_805;
      end
      11'b01100100110 : begin
        result = input_806;
      end
      11'b01100100111 : begin
        result = input_807;
      end
      11'b01100101000 : begin
        result = input_808;
      end
      11'b01100101001 : begin
        result = input_809;
      end
      11'b01100101010 : begin
        result = input_810;
      end
      11'b01100101011 : begin
        result = input_811;
      end
      11'b01100101100 : begin
        result = input_812;
      end
      11'b01100101101 : begin
        result = input_813;
      end
      11'b01100101110 : begin
        result = input_814;
      end
      11'b01100101111 : begin
        result = input_815;
      end
      11'b01100110000 : begin
        result = input_816;
      end
      11'b01100110001 : begin
        result = input_817;
      end
      11'b01100110010 : begin
        result = input_818;
      end
      11'b01100110011 : begin
        result = input_819;
      end
      11'b01100110100 : begin
        result = input_820;
      end
      11'b01100110101 : begin
        result = input_821;
      end
      11'b01100110110 : begin
        result = input_822;
      end
      11'b01100110111 : begin
        result = input_823;
      end
      11'b01100111000 : begin
        result = input_824;
      end
      11'b01100111001 : begin
        result = input_825;
      end
      11'b01100111010 : begin
        result = input_826;
      end
      11'b01100111011 : begin
        result = input_827;
      end
      11'b01100111100 : begin
        result = input_828;
      end
      11'b01100111101 : begin
        result = input_829;
      end
      11'b01100111110 : begin
        result = input_830;
      end
      11'b01100111111 : begin
        result = input_831;
      end
      11'b01101000000 : begin
        result = input_832;
      end
      11'b01101000001 : begin
        result = input_833;
      end
      11'b01101000010 : begin
        result = input_834;
      end
      11'b01101000011 : begin
        result = input_835;
      end
      11'b01101000100 : begin
        result = input_836;
      end
      11'b01101000101 : begin
        result = input_837;
      end
      11'b01101000110 : begin
        result = input_838;
      end
      11'b01101000111 : begin
        result = input_839;
      end
      11'b01101001000 : begin
        result = input_840;
      end
      11'b01101001001 : begin
        result = input_841;
      end
      11'b01101001010 : begin
        result = input_842;
      end
      11'b01101001011 : begin
        result = input_843;
      end
      11'b01101001100 : begin
        result = input_844;
      end
      11'b01101001101 : begin
        result = input_845;
      end
      11'b01101001110 : begin
        result = input_846;
      end
      11'b01101001111 : begin
        result = input_847;
      end
      11'b01101010000 : begin
        result = input_848;
      end
      11'b01101010001 : begin
        result = input_849;
      end
      11'b01101010010 : begin
        result = input_850;
      end
      11'b01101010011 : begin
        result = input_851;
      end
      11'b01101010100 : begin
        result = input_852;
      end
      11'b01101010101 : begin
        result = input_853;
      end
      11'b01101010110 : begin
        result = input_854;
      end
      11'b01101010111 : begin
        result = input_855;
      end
      11'b01101011000 : begin
        result = input_856;
      end
      11'b01101011001 : begin
        result = input_857;
      end
      11'b01101011010 : begin
        result = input_858;
      end
      11'b01101011011 : begin
        result = input_859;
      end
      11'b01101011100 : begin
        result = input_860;
      end
      11'b01101011101 : begin
        result = input_861;
      end
      11'b01101011110 : begin
        result = input_862;
      end
      11'b01101011111 : begin
        result = input_863;
      end
      11'b01101100000 : begin
        result = input_864;
      end
      11'b01101100001 : begin
        result = input_865;
      end
      11'b01101100010 : begin
        result = input_866;
      end
      11'b01101100011 : begin
        result = input_867;
      end
      11'b01101100100 : begin
        result = input_868;
      end
      11'b01101100101 : begin
        result = input_869;
      end
      11'b01101100110 : begin
        result = input_870;
      end
      11'b01101100111 : begin
        result = input_871;
      end
      11'b01101101000 : begin
        result = input_872;
      end
      11'b01101101001 : begin
        result = input_873;
      end
      11'b01101101010 : begin
        result = input_874;
      end
      11'b01101101011 : begin
        result = input_875;
      end
      11'b01101101100 : begin
        result = input_876;
      end
      11'b01101101101 : begin
        result = input_877;
      end
      11'b01101101110 : begin
        result = input_878;
      end
      11'b01101101111 : begin
        result = input_879;
      end
      11'b01101110000 : begin
        result = input_880;
      end
      11'b01101110001 : begin
        result = input_881;
      end
      11'b01101110010 : begin
        result = input_882;
      end
      11'b01101110011 : begin
        result = input_883;
      end
      11'b01101110100 : begin
        result = input_884;
      end
      11'b01101110101 : begin
        result = input_885;
      end
      11'b01101110110 : begin
        result = input_886;
      end
      11'b01101110111 : begin
        result = input_887;
      end
      11'b01101111000 : begin
        result = input_888;
      end
      11'b01101111001 : begin
        result = input_889;
      end
      11'b01101111010 : begin
        result = input_890;
      end
      11'b01101111011 : begin
        result = input_891;
      end
      11'b01101111100 : begin
        result = input_892;
      end
      11'b01101111101 : begin
        result = input_893;
      end
      11'b01101111110 : begin
        result = input_894;
      end
      11'b01101111111 : begin
        result = input_895;
      end
      11'b01110000000 : begin
        result = input_896;
      end
      11'b01110000001 : begin
        result = input_897;
      end
      11'b01110000010 : begin
        result = input_898;
      end
      11'b01110000011 : begin
        result = input_899;
      end
      11'b01110000100 : begin
        result = input_900;
      end
      11'b01110000101 : begin
        result = input_901;
      end
      11'b01110000110 : begin
        result = input_902;
      end
      11'b01110000111 : begin
        result = input_903;
      end
      11'b01110001000 : begin
        result = input_904;
      end
      11'b01110001001 : begin
        result = input_905;
      end
      11'b01110001010 : begin
        result = input_906;
      end
      11'b01110001011 : begin
        result = input_907;
      end
      11'b01110001100 : begin
        result = input_908;
      end
      11'b01110001101 : begin
        result = input_909;
      end
      11'b01110001110 : begin
        result = input_910;
      end
      11'b01110001111 : begin
        result = input_911;
      end
      11'b01110010000 : begin
        result = input_912;
      end
      11'b01110010001 : begin
        result = input_913;
      end
      11'b01110010010 : begin
        result = input_914;
      end
      11'b01110010011 : begin
        result = input_915;
      end
      11'b01110010100 : begin
        result = input_916;
      end
      11'b01110010101 : begin
        result = input_917;
      end
      11'b01110010110 : begin
        result = input_918;
      end
      11'b01110010111 : begin
        result = input_919;
      end
      11'b01110011000 : begin
        result = input_920;
      end
      11'b01110011001 : begin
        result = input_921;
      end
      11'b01110011010 : begin
        result = input_922;
      end
      11'b01110011011 : begin
        result = input_923;
      end
      11'b01110011100 : begin
        result = input_924;
      end
      11'b01110011101 : begin
        result = input_925;
      end
      11'b01110011110 : begin
        result = input_926;
      end
      11'b01110011111 : begin
        result = input_927;
      end
      11'b01110100000 : begin
        result = input_928;
      end
      11'b01110100001 : begin
        result = input_929;
      end
      11'b01110100010 : begin
        result = input_930;
      end
      11'b01110100011 : begin
        result = input_931;
      end
      11'b01110100100 : begin
        result = input_932;
      end
      11'b01110100101 : begin
        result = input_933;
      end
      11'b01110100110 : begin
        result = input_934;
      end
      11'b01110100111 : begin
        result = input_935;
      end
      11'b01110101000 : begin
        result = input_936;
      end
      11'b01110101001 : begin
        result = input_937;
      end
      11'b01110101010 : begin
        result = input_938;
      end
      11'b01110101011 : begin
        result = input_939;
      end
      11'b01110101100 : begin
        result = input_940;
      end
      11'b01110101101 : begin
        result = input_941;
      end
      11'b01110101110 : begin
        result = input_942;
      end
      11'b01110101111 : begin
        result = input_943;
      end
      11'b01110110000 : begin
        result = input_944;
      end
      11'b01110110001 : begin
        result = input_945;
      end
      11'b01110110010 : begin
        result = input_946;
      end
      11'b01110110011 : begin
        result = input_947;
      end
      11'b01110110100 : begin
        result = input_948;
      end
      11'b01110110101 : begin
        result = input_949;
      end
      11'b01110110110 : begin
        result = input_950;
      end
      11'b01110110111 : begin
        result = input_951;
      end
      11'b01110111000 : begin
        result = input_952;
      end
      11'b01110111001 : begin
        result = input_953;
      end
      11'b01110111010 : begin
        result = input_954;
      end
      11'b01110111011 : begin
        result = input_955;
      end
      11'b01110111100 : begin
        result = input_956;
      end
      11'b01110111101 : begin
        result = input_957;
      end
      11'b01110111110 : begin
        result = input_958;
      end
      11'b01110111111 : begin
        result = input_959;
      end
      11'b01111000000 : begin
        result = input_960;
      end
      11'b01111000001 : begin
        result = input_961;
      end
      11'b01111000010 : begin
        result = input_962;
      end
      11'b01111000011 : begin
        result = input_963;
      end
      11'b01111000100 : begin
        result = input_964;
      end
      11'b01111000101 : begin
        result = input_965;
      end
      11'b01111000110 : begin
        result = input_966;
      end
      11'b01111000111 : begin
        result = input_967;
      end
      11'b01111001000 : begin
        result = input_968;
      end
      11'b01111001001 : begin
        result = input_969;
      end
      11'b01111001010 : begin
        result = input_970;
      end
      11'b01111001011 : begin
        result = input_971;
      end
      11'b01111001100 : begin
        result = input_972;
      end
      11'b01111001101 : begin
        result = input_973;
      end
      11'b01111001110 : begin
        result = input_974;
      end
      11'b01111001111 : begin
        result = input_975;
      end
      11'b01111010000 : begin
        result = input_976;
      end
      11'b01111010001 : begin
        result = input_977;
      end
      11'b01111010010 : begin
        result = input_978;
      end
      11'b01111010011 : begin
        result = input_979;
      end
      11'b01111010100 : begin
        result = input_980;
      end
      11'b01111010101 : begin
        result = input_981;
      end
      11'b01111010110 : begin
        result = input_982;
      end
      11'b01111010111 : begin
        result = input_983;
      end
      11'b01111011000 : begin
        result = input_984;
      end
      11'b01111011001 : begin
        result = input_985;
      end
      11'b01111011010 : begin
        result = input_986;
      end
      11'b01111011011 : begin
        result = input_987;
      end
      11'b01111011100 : begin
        result = input_988;
      end
      11'b01111011101 : begin
        result = input_989;
      end
      11'b01111011110 : begin
        result = input_990;
      end
      11'b01111011111 : begin
        result = input_991;
      end
      11'b01111100000 : begin
        result = input_992;
      end
      11'b01111100001 : begin
        result = input_993;
      end
      11'b01111100010 : begin
        result = input_994;
      end
      11'b01111100011 : begin
        result = input_995;
      end
      11'b01111100100 : begin
        result = input_996;
      end
      11'b01111100101 : begin
        result = input_997;
      end
      11'b01111100110 : begin
        result = input_998;
      end
      11'b01111100111 : begin
        result = input_999;
      end
      11'b01111101000 : begin
        result = input_1000;
      end
      11'b01111101001 : begin
        result = input_1001;
      end
      11'b01111101010 : begin
        result = input_1002;
      end
      11'b01111101011 : begin
        result = input_1003;
      end
      11'b01111101100 : begin
        result = input_1004;
      end
      11'b01111101101 : begin
        result = input_1005;
      end
      11'b01111101110 : begin
        result = input_1006;
      end
      11'b01111101111 : begin
        result = input_1007;
      end
      11'b01111110000 : begin
        result = input_1008;
      end
      11'b01111110001 : begin
        result = input_1009;
      end
      11'b01111110010 : begin
        result = input_1010;
      end
      11'b01111110011 : begin
        result = input_1011;
      end
      11'b01111110100 : begin
        result = input_1012;
      end
      11'b01111110101 : begin
        result = input_1013;
      end
      11'b01111110110 : begin
        result = input_1014;
      end
      11'b01111110111 : begin
        result = input_1015;
      end
      11'b01111111000 : begin
        result = input_1016;
      end
      11'b01111111001 : begin
        result = input_1017;
      end
      11'b01111111010 : begin
        result = input_1018;
      end
      11'b01111111011 : begin
        result = input_1019;
      end
      11'b01111111100 : begin
        result = input_1020;
      end
      11'b01111111101 : begin
        result = input_1021;
      end
      11'b01111111110 : begin
        result = input_1022;
      end
      11'b01111111111 : begin
        result = input_1023;
      end
      11'b10000000000 : begin
        result = input_1024;
      end
      11'b10000000001 : begin
        result = input_1025;
      end
      11'b10000000010 : begin
        result = input_1026;
      end
      11'b10000000011 : begin
        result = input_1027;
      end
      11'b10000000100 : begin
        result = input_1028;
      end
      11'b10000000101 : begin
        result = input_1029;
      end
      11'b10000000110 : begin
        result = input_1030;
      end
      11'b10000000111 : begin
        result = input_1031;
      end
      11'b10000001000 : begin
        result = input_1032;
      end
      11'b10000001001 : begin
        result = input_1033;
      end
      11'b10000001010 : begin
        result = input_1034;
      end
      11'b10000001011 : begin
        result = input_1035;
      end
      11'b10000001100 : begin
        result = input_1036;
      end
      11'b10000001101 : begin
        result = input_1037;
      end
      11'b10000001110 : begin
        result = input_1038;
      end
      11'b10000001111 : begin
        result = input_1039;
      end
      11'b10000010000 : begin
        result = input_1040;
      end
      11'b10000010001 : begin
        result = input_1041;
      end
      11'b10000010010 : begin
        result = input_1042;
      end
      11'b10000010011 : begin
        result = input_1043;
      end
      11'b10000010100 : begin
        result = input_1044;
      end
      11'b10000010101 : begin
        result = input_1045;
      end
      11'b10000010110 : begin
        result = input_1046;
      end
      11'b10000010111 : begin
        result = input_1047;
      end
      11'b10000011000 : begin
        result = input_1048;
      end
      11'b10000011001 : begin
        result = input_1049;
      end
      11'b10000011010 : begin
        result = input_1050;
      end
      11'b10000011011 : begin
        result = input_1051;
      end
      11'b10000011100 : begin
        result = input_1052;
      end
      11'b10000011101 : begin
        result = input_1053;
      end
      11'b10000011110 : begin
        result = input_1054;
      end
      11'b10000011111 : begin
        result = input_1055;
      end
      11'b10000100000 : begin
        result = input_1056;
      end
      11'b10000100001 : begin
        result = input_1057;
      end
      11'b10000100010 : begin
        result = input_1058;
      end
      11'b10000100011 : begin
        result = input_1059;
      end
      11'b10000100100 : begin
        result = input_1060;
      end
      11'b10000100101 : begin
        result = input_1061;
      end
      11'b10000100110 : begin
        result = input_1062;
      end
      11'b10000100111 : begin
        result = input_1063;
      end
      11'b10000101000 : begin
        result = input_1064;
      end
      11'b10000101001 : begin
        result = input_1065;
      end
      11'b10000101010 : begin
        result = input_1066;
      end
      11'b10000101011 : begin
        result = input_1067;
      end
      11'b10000101100 : begin
        result = input_1068;
      end
      11'b10000101101 : begin
        result = input_1069;
      end
      11'b10000101110 : begin
        result = input_1070;
      end
      11'b10000101111 : begin
        result = input_1071;
      end
      11'b10000110000 : begin
        result = input_1072;
      end
      11'b10000110001 : begin
        result = input_1073;
      end
      11'b10000110010 : begin
        result = input_1074;
      end
      11'b10000110011 : begin
        result = input_1075;
      end
      11'b10000110100 : begin
        result = input_1076;
      end
      11'b10000110101 : begin
        result = input_1077;
      end
      11'b10000110110 : begin
        result = input_1078;
      end
      11'b10000110111 : begin
        result = input_1079;
      end
      11'b10000111000 : begin
        result = input_1080;
      end
      11'b10000111001 : begin
        result = input_1081;
      end
      11'b10000111010 : begin
        result = input_1082;
      end
      11'b10000111011 : begin
        result = input_1083;
      end
      11'b10000111100 : begin
        result = input_1084;
      end
      11'b10000111101 : begin
        result = input_1085;
      end
      11'b10000111110 : begin
        result = input_1086;
      end
      11'b10000111111 : begin
        result = input_1087;
      end
      11'b10001000000 : begin
        result = input_1088;
      end
      11'b10001000001 : begin
        result = input_1089;
      end
      11'b10001000010 : begin
        result = input_1090;
      end
      11'b10001000011 : begin
        result = input_1091;
      end
      11'b10001000100 : begin
        result = input_1092;
      end
      11'b10001000101 : begin
        result = input_1093;
      end
      11'b10001000110 : begin
        result = input_1094;
      end
      11'b10001000111 : begin
        result = input_1095;
      end
      11'b10001001000 : begin
        result = input_1096;
      end
      11'b10001001001 : begin
        result = input_1097;
      end
      11'b10001001010 : begin
        result = input_1098;
      end
      11'b10001001011 : begin
        result = input_1099;
      end
      11'b10001001100 : begin
        result = input_1100;
      end
      11'b10001001101 : begin
        result = input_1101;
      end
      11'b10001001110 : begin
        result = input_1102;
      end
      11'b10001001111 : begin
        result = input_1103;
      end
      11'b10001010000 : begin
        result = input_1104;
      end
      11'b10001010001 : begin
        result = input_1105;
      end
      11'b10001010010 : begin
        result = input_1106;
      end
      11'b10001010011 : begin
        result = input_1107;
      end
      11'b10001010100 : begin
        result = input_1108;
      end
      11'b10001010101 : begin
        result = input_1109;
      end
      11'b10001010110 : begin
        result = input_1110;
      end
      11'b10001010111 : begin
        result = input_1111;
      end
      11'b10001011000 : begin
        result = input_1112;
      end
      11'b10001011001 : begin
        result = input_1113;
      end
      11'b10001011010 : begin
        result = input_1114;
      end
      11'b10001011011 : begin
        result = input_1115;
      end
      11'b10001011100 : begin
        result = input_1116;
      end
      11'b10001011101 : begin
        result = input_1117;
      end
      11'b10001011110 : begin
        result = input_1118;
      end
      11'b10001011111 : begin
        result = input_1119;
      end
      11'b10001100000 : begin
        result = input_1120;
      end
      11'b10001100001 : begin
        result = input_1121;
      end
      11'b10001100010 : begin
        result = input_1122;
      end
      11'b10001100011 : begin
        result = input_1123;
      end
      11'b10001100100 : begin
        result = input_1124;
      end
      11'b10001100101 : begin
        result = input_1125;
      end
      11'b10001100110 : begin
        result = input_1126;
      end
      11'b10001100111 : begin
        result = input_1127;
      end
      11'b10001101000 : begin
        result = input_1128;
      end
      11'b10001101001 : begin
        result = input_1129;
      end
      11'b10001101010 : begin
        result = input_1130;
      end
      11'b10001101011 : begin
        result = input_1131;
      end
      11'b10001101100 : begin
        result = input_1132;
      end
      11'b10001101101 : begin
        result = input_1133;
      end
      11'b10001101110 : begin
        result = input_1134;
      end
      11'b10001101111 : begin
        result = input_1135;
      end
      11'b10001110000 : begin
        result = input_1136;
      end
      11'b10001110001 : begin
        result = input_1137;
      end
      11'b10001110010 : begin
        result = input_1138;
      end
      11'b10001110011 : begin
        result = input_1139;
      end
      11'b10001110100 : begin
        result = input_1140;
      end
      11'b10001110101 : begin
        result = input_1141;
      end
      11'b10001110110 : begin
        result = input_1142;
      end
      11'b10001110111 : begin
        result = input_1143;
      end
      11'b10001111000 : begin
        result = input_1144;
      end
      11'b10001111001 : begin
        result = input_1145;
      end
      11'b10001111010 : begin
        result = input_1146;
      end
      11'b10001111011 : begin
        result = input_1147;
      end
      11'b10001111100 : begin
        result = input_1148;
      end
      11'b10001111101 : begin
        result = input_1149;
      end
      11'b10001111110 : begin
        result = input_1150;
      end
      11'b10001111111 : begin
        result = input_1151;
      end
      11'b10010000000 : begin
        result = input_1152;
      end
      11'b10010000001 : begin
        result = input_1153;
      end
      11'b10010000010 : begin
        result = input_1154;
      end
      11'b10010000011 : begin
        result = input_1155;
      end
      11'b10010000100 : begin
        result = input_1156;
      end
      11'b10010000101 : begin
        result = input_1157;
      end
      11'b10010000110 : begin
        result = input_1158;
      end
      11'b10010000111 : begin
        result = input_1159;
      end
      11'b10010001000 : begin
        result = input_1160;
      end
      11'b10010001001 : begin
        result = input_1161;
      end
      11'b10010001010 : begin
        result = input_1162;
      end
      11'b10010001011 : begin
        result = input_1163;
      end
      11'b10010001100 : begin
        result = input_1164;
      end
      11'b10010001101 : begin
        result = input_1165;
      end
      11'b10010001110 : begin
        result = input_1166;
      end
      11'b10010001111 : begin
        result = input_1167;
      end
      11'b10010010000 : begin
        result = input_1168;
      end
      11'b10010010001 : begin
        result = input_1169;
      end
      11'b10010010010 : begin
        result = input_1170;
      end
      11'b10010010011 : begin
        result = input_1171;
      end
      11'b10010010100 : begin
        result = input_1172;
      end
      11'b10010010101 : begin
        result = input_1173;
      end
      11'b10010010110 : begin
        result = input_1174;
      end
      11'b10010010111 : begin
        result = input_1175;
      end
      11'b10010011000 : begin
        result = input_1176;
      end
      11'b10010011001 : begin
        result = input_1177;
      end
      11'b10010011010 : begin
        result = input_1178;
      end
      11'b10010011011 : begin
        result = input_1179;
      end
      11'b10010011100 : begin
        result = input_1180;
      end
      11'b10010011101 : begin
        result = input_1181;
      end
      11'b10010011110 : begin
        result = input_1182;
      end
      11'b10010011111 : begin
        result = input_1183;
      end
      11'b10010100000 : begin
        result = input_1184;
      end
      11'b10010100001 : begin
        result = input_1185;
      end
      11'b10010100010 : begin
        result = input_1186;
      end
      11'b10010100011 : begin
        result = input_1187;
      end
      11'b10010100100 : begin
        result = input_1188;
      end
      11'b10010100101 : begin
        result = input_1189;
      end
      11'b10010100110 : begin
        result = input_1190;
      end
      11'b10010100111 : begin
        result = input_1191;
      end
      11'b10010101000 : begin
        result = input_1192;
      end
      11'b10010101001 : begin
        result = input_1193;
      end
      11'b10010101010 : begin
        result = input_1194;
      end
      11'b10010101011 : begin
        result = input_1195;
      end
      11'b10010101100 : begin
        result = input_1196;
      end
      11'b10010101101 : begin
        result = input_1197;
      end
      11'b10010101110 : begin
        result = input_1198;
      end
      11'b10010101111 : begin
        result = input_1199;
      end
      11'b10010110000 : begin
        result = input_1200;
      end
      11'b10010110001 : begin
        result = input_1201;
      end
      11'b10010110010 : begin
        result = input_1202;
      end
      11'b10010110011 : begin
        result = input_1203;
      end
      11'b10010110100 : begin
        result = input_1204;
      end
      11'b10010110101 : begin
        result = input_1205;
      end
      11'b10010110110 : begin
        result = input_1206;
      end
      11'b10010110111 : begin
        result = input_1207;
      end
      11'b10010111000 : begin
        result = input_1208;
      end
      11'b10010111001 : begin
        result = input_1209;
      end
      11'b10010111010 : begin
        result = input_1210;
      end
      11'b10010111011 : begin
        result = input_1211;
      end
      11'b10010111100 : begin
        result = input_1212;
      end
      11'b10010111101 : begin
        result = input_1213;
      end
      11'b10010111110 : begin
        result = input_1214;
      end
      11'b10010111111 : begin
        result = input_1215;
      end
      11'b10011000000 : begin
        result = input_1216;
      end
      11'b10011000001 : begin
        result = input_1217;
      end
      11'b10011000010 : begin
        result = input_1218;
      end
      11'b10011000011 : begin
        result = input_1219;
      end
      11'b10011000100 : begin
        result = input_1220;
      end
      11'b10011000101 : begin
        result = input_1221;
      end
      11'b10011000110 : begin
        result = input_1222;
      end
      11'b10011000111 : begin
        result = input_1223;
      end
      11'b10011001000 : begin
        result = input_1224;
      end
      11'b10011001001 : begin
        result = input_1225;
      end
      11'b10011001010 : begin
        result = input_1226;
      end
      11'b10011001011 : begin
        result = input_1227;
      end
      11'b10011001100 : begin
        result = input_1228;
      end
      11'b10011001101 : begin
        result = input_1229;
      end
      11'b10011001110 : begin
        result = input_1230;
      end
      11'b10011001111 : begin
        result = input_1231;
      end
      11'b10011010000 : begin
        result = input_1232;
      end
      11'b10011010001 : begin
        result = input_1233;
      end
      11'b10011010010 : begin
        result = input_1234;
      end
      11'b10011010011 : begin
        result = input_1235;
      end
      11'b10011010100 : begin
        result = input_1236;
      end
      11'b10011010101 : begin
        result = input_1237;
      end
      11'b10011010110 : begin
        result = input_1238;
      end
      11'b10011010111 : begin
        result = input_1239;
      end
      11'b10011011000 : begin
        result = input_1240;
      end
      11'b10011011001 : begin
        result = input_1241;
      end
      11'b10011011010 : begin
        result = input_1242;
      end
      11'b10011011011 : begin
        result = input_1243;
      end
      11'b10011011100 : begin
        result = input_1244;
      end
      11'b10011011101 : begin
        result = input_1245;
      end
      11'b10011011110 : begin
        result = input_1246;
      end
      11'b10011011111 : begin
        result = input_1247;
      end
      11'b10011100000 : begin
        result = input_1248;
      end
      11'b10011100001 : begin
        result = input_1249;
      end
      11'b10011100010 : begin
        result = input_1250;
      end
      11'b10011100011 : begin
        result = input_1251;
      end
      11'b10011100100 : begin
        result = input_1252;
      end
      11'b10011100101 : begin
        result = input_1253;
      end
      11'b10011100110 : begin
        result = input_1254;
      end
      11'b10011100111 : begin
        result = input_1255;
      end
      11'b10011101000 : begin
        result = input_1256;
      end
      11'b10011101001 : begin
        result = input_1257;
      end
      11'b10011101010 : begin
        result = input_1258;
      end
      11'b10011101011 : begin
        result = input_1259;
      end
      11'b10011101100 : begin
        result = input_1260;
      end
      11'b10011101101 : begin
        result = input_1261;
      end
      11'b10011101110 : begin
        result = input_1262;
      end
      11'b10011101111 : begin
        result = input_1263;
      end
      11'b10011110000 : begin
        result = input_1264;
      end
      11'b10011110001 : begin
        result = input_1265;
      end
      11'b10011110010 : begin
        result = input_1266;
      end
      11'b10011110011 : begin
        result = input_1267;
      end
      11'b10011110100 : begin
        result = input_1268;
      end
      11'b10011110101 : begin
        result = input_1269;
      end
      11'b10011110110 : begin
        result = input_1270;
      end
      11'b10011110111 : begin
        result = input_1271;
      end
      11'b10011111000 : begin
        result = input_1272;
      end
      11'b10011111001 : begin
        result = input_1273;
      end
      11'b10011111010 : begin
        result = input_1274;
      end
      11'b10011111011 : begin
        result = input_1275;
      end
      11'b10011111100 : begin
        result = input_1276;
      end
      11'b10011111101 : begin
        result = input_1277;
      end
      11'b10011111110 : begin
        result = input_1278;
      end
      11'b10011111111 : begin
        result = input_1279;
      end
      11'b10100000000 : begin
        result = input_1280;
      end
      11'b10100000001 : begin
        result = input_1281;
      end
      11'b10100000010 : begin
        result = input_1282;
      end
      11'b10100000011 : begin
        result = input_1283;
      end
      11'b10100000100 : begin
        result = input_1284;
      end
      11'b10100000101 : begin
        result = input_1285;
      end
      11'b10100000110 : begin
        result = input_1286;
      end
      11'b10100000111 : begin
        result = input_1287;
      end
      11'b10100001000 : begin
        result = input_1288;
      end
      11'b10100001001 : begin
        result = input_1289;
      end
      11'b10100001010 : begin
        result = input_1290;
      end
      11'b10100001011 : begin
        result = input_1291;
      end
      11'b10100001100 : begin
        result = input_1292;
      end
      11'b10100001101 : begin
        result = input_1293;
      end
      11'b10100001110 : begin
        result = input_1294;
      end
      11'b10100001111 : begin
        result = input_1295;
      end
      11'b10100010000 : begin
        result = input_1296;
      end
      11'b10100010001 : begin
        result = input_1297;
      end
      11'b10100010010 : begin
        result = input_1298;
      end
      11'b10100010011 : begin
        result = input_1299;
      end
      11'b10100010100 : begin
        result = input_1300;
      end
      11'b10100010101 : begin
        result = input_1301;
      end
      11'b10100010110 : begin
        result = input_1302;
      end
      11'b10100010111 : begin
        result = input_1303;
      end
      11'b10100011000 : begin
        result = input_1304;
      end
      11'b10100011001 : begin
        result = input_1305;
      end
      11'b10100011010 : begin
        result = input_1306;
      end
      11'b10100011011 : begin
        result = input_1307;
      end
      11'b10100011100 : begin
        result = input_1308;
      end
      11'b10100011101 : begin
        result = input_1309;
      end
      11'b10100011110 : begin
        result = input_1310;
      end
      11'b10100011111 : begin
        result = input_1311;
      end
      11'b10100100000 : begin
        result = input_1312;
      end
      11'b10100100001 : begin
        result = input_1313;
      end
      11'b10100100010 : begin
        result = input_1314;
      end
      11'b10100100011 : begin
        result = input_1315;
      end
      11'b10100100100 : begin
        result = input_1316;
      end
      11'b10100100101 : begin
        result = input_1317;
      end
      11'b10100100110 : begin
        result = input_1318;
      end
      11'b10100100111 : begin
        result = input_1319;
      end
      11'b10100101000 : begin
        result = input_1320;
      end
      11'b10100101001 : begin
        result = input_1321;
      end
      11'b10100101010 : begin
        result = input_1322;
      end
      11'b10100101011 : begin
        result = input_1323;
      end
      11'b10100101100 : begin
        result = input_1324;
      end
      11'b10100101101 : begin
        result = input_1325;
      end
      11'b10100101110 : begin
        result = input_1326;
      end
      11'b10100101111 : begin
        result = input_1327;
      end
      11'b10100110000 : begin
        result = input_1328;
      end
      11'b10100110001 : begin
        result = input_1329;
      end
      11'b10100110010 : begin
        result = input_1330;
      end
      11'b10100110011 : begin
        result = input_1331;
      end
      11'b10100110100 : begin
        result = input_1332;
      end
      11'b10100110101 : begin
        result = input_1333;
      end
      11'b10100110110 : begin
        result = input_1334;
      end
      11'b10100110111 : begin
        result = input_1335;
      end
      11'b10100111000 : begin
        result = input_1336;
      end
      11'b10100111001 : begin
        result = input_1337;
      end
      11'b10100111010 : begin
        result = input_1338;
      end
      11'b10100111011 : begin
        result = input_1339;
      end
      11'b10100111100 : begin
        result = input_1340;
      end
      11'b10100111101 : begin
        result = input_1341;
      end
      11'b10100111110 : begin
        result = input_1342;
      end
      11'b10100111111 : begin
        result = input_1343;
      end
      11'b10101000000 : begin
        result = input_1344;
      end
      11'b10101000001 : begin
        result = input_1345;
      end
      11'b10101000010 : begin
        result = input_1346;
      end
      11'b10101000011 : begin
        result = input_1347;
      end
      11'b10101000100 : begin
        result = input_1348;
      end
      11'b10101000101 : begin
        result = input_1349;
      end
      11'b10101000110 : begin
        result = input_1350;
      end
      11'b10101000111 : begin
        result = input_1351;
      end
      11'b10101001000 : begin
        result = input_1352;
      end
      11'b10101001001 : begin
        result = input_1353;
      end
      11'b10101001010 : begin
        result = input_1354;
      end
      11'b10101001011 : begin
        result = input_1355;
      end
      11'b10101001100 : begin
        result = input_1356;
      end
      11'b10101001101 : begin
        result = input_1357;
      end
      11'b10101001110 : begin
        result = input_1358;
      end
      11'b10101001111 : begin
        result = input_1359;
      end
      11'b10101010000 : begin
        result = input_1360;
      end
      11'b10101010001 : begin
        result = input_1361;
      end
      11'b10101010010 : begin
        result = input_1362;
      end
      11'b10101010011 : begin
        result = input_1363;
      end
      11'b10101010100 : begin
        result = input_1364;
      end
      11'b10101010101 : begin
        result = input_1365;
      end
      11'b10101010110 : begin
        result = input_1366;
      end
      11'b10101010111 : begin
        result = input_1367;
      end
      11'b10101011000 : begin
        result = input_1368;
      end
      11'b10101011001 : begin
        result = input_1369;
      end
      11'b10101011010 : begin
        result = input_1370;
      end
      11'b10101011011 : begin
        result = input_1371;
      end
      11'b10101011100 : begin
        result = input_1372;
      end
      11'b10101011101 : begin
        result = input_1373;
      end
      11'b10101011110 : begin
        result = input_1374;
      end
      11'b10101011111 : begin
        result = input_1375;
      end
      11'b10101100000 : begin
        result = input_1376;
      end
      11'b10101100001 : begin
        result = input_1377;
      end
      11'b10101100010 : begin
        result = input_1378;
      end
      11'b10101100011 : begin
        result = input_1379;
      end
      11'b10101100100 : begin
        result = input_1380;
      end
      11'b10101100101 : begin
        result = input_1381;
      end
      11'b10101100110 : begin
        result = input_1382;
      end
      11'b10101100111 : begin
        result = input_1383;
      end
      11'b10101101000 : begin
        result = input_1384;
      end
      11'b10101101001 : begin
        result = input_1385;
      end
      11'b10101101010 : begin
        result = input_1386;
      end
      11'b10101101011 : begin
        result = input_1387;
      end
      11'b10101101100 : begin
        result = input_1388;
      end
      11'b10101101101 : begin
        result = input_1389;
      end
      11'b10101101110 : begin
        result = input_1390;
      end
      11'b10101101111 : begin
        result = input_1391;
      end
      11'b10101110000 : begin
        result = input_1392;
      end
      11'b10101110001 : begin
        result = input_1393;
      end
      11'b10101110010 : begin
        result = input_1394;
      end
      11'b10101110011 : begin
        result = input_1395;
      end
      11'b10101110100 : begin
        result = input_1396;
      end
      11'b10101110101 : begin
        result = input_1397;
      end
      11'b10101110110 : begin
        result = input_1398;
      end
      11'b10101110111 : begin
        result = input_1399;
      end
      11'b10101111000 : begin
        result = input_1400;
      end
      11'b10101111001 : begin
        result = input_1401;
      end
      11'b10101111010 : begin
        result = input_1402;
      end
      11'b10101111011 : begin
        result = input_1403;
      end
      11'b10101111100 : begin
        result = input_1404;
      end
      11'b10101111101 : begin
        result = input_1405;
      end
      11'b10101111110 : begin
        result = input_1406;
      end
      11'b10101111111 : begin
        result = input_1407;
      end
      11'b10110000000 : begin
        result = input_1408;
      end
      11'b10110000001 : begin
        result = input_1409;
      end
      11'b10110000010 : begin
        result = input_1410;
      end
      11'b10110000011 : begin
        result = input_1411;
      end
      11'b10110000100 : begin
        result = input_1412;
      end
      11'b10110000101 : begin
        result = input_1413;
      end
      11'b10110000110 : begin
        result = input_1414;
      end
      11'b10110000111 : begin
        result = input_1415;
      end
      11'b10110001000 : begin
        result = input_1416;
      end
      11'b10110001001 : begin
        result = input_1417;
      end
      11'b10110001010 : begin
        result = input_1418;
      end
      11'b10110001011 : begin
        result = input_1419;
      end
      11'b10110001100 : begin
        result = input_1420;
      end
      11'b10110001101 : begin
        result = input_1421;
      end
      11'b10110001110 : begin
        result = input_1422;
      end
      11'b10110001111 : begin
        result = input_1423;
      end
      11'b10110010000 : begin
        result = input_1424;
      end
      11'b10110010001 : begin
        result = input_1425;
      end
      11'b10110010010 : begin
        result = input_1426;
      end
      11'b10110010011 : begin
        result = input_1427;
      end
      11'b10110010100 : begin
        result = input_1428;
      end
      11'b10110010101 : begin
        result = input_1429;
      end
      11'b10110010110 : begin
        result = input_1430;
      end
      11'b10110010111 : begin
        result = input_1431;
      end
      11'b10110011000 : begin
        result = input_1432;
      end
      11'b10110011001 : begin
        result = input_1433;
      end
      11'b10110011010 : begin
        result = input_1434;
      end
      11'b10110011011 : begin
        result = input_1435;
      end
      11'b10110011100 : begin
        result = input_1436;
      end
      11'b10110011101 : begin
        result = input_1437;
      end
      11'b10110011110 : begin
        result = input_1438;
      end
      11'b10110011111 : begin
        result = input_1439;
      end
      11'b10110100000 : begin
        result = input_1440;
      end
      11'b10110100001 : begin
        result = input_1441;
      end
      11'b10110100010 : begin
        result = input_1442;
      end
      11'b10110100011 : begin
        result = input_1443;
      end
      11'b10110100100 : begin
        result = input_1444;
      end
      11'b10110100101 : begin
        result = input_1445;
      end
      11'b10110100110 : begin
        result = input_1446;
      end
      11'b10110100111 : begin
        result = input_1447;
      end
      11'b10110101000 : begin
        result = input_1448;
      end
      11'b10110101001 : begin
        result = input_1449;
      end
      11'b10110101010 : begin
        result = input_1450;
      end
      11'b10110101011 : begin
        result = input_1451;
      end
      11'b10110101100 : begin
        result = input_1452;
      end
      11'b10110101101 : begin
        result = input_1453;
      end
      11'b10110101110 : begin
        result = input_1454;
      end
      11'b10110101111 : begin
        result = input_1455;
      end
      11'b10110110000 : begin
        result = input_1456;
      end
      11'b10110110001 : begin
        result = input_1457;
      end
      11'b10110110010 : begin
        result = input_1458;
      end
      11'b10110110011 : begin
        result = input_1459;
      end
      11'b10110110100 : begin
        result = input_1460;
      end
      11'b10110110101 : begin
        result = input_1461;
      end
      11'b10110110110 : begin
        result = input_1462;
      end
      11'b10110110111 : begin
        result = input_1463;
      end
      11'b10110111000 : begin
        result = input_1464;
      end
      11'b10110111001 : begin
        result = input_1465;
      end
      11'b10110111010 : begin
        result = input_1466;
      end
      11'b10110111011 : begin
        result = input_1467;
      end
      11'b10110111100 : begin
        result = input_1468;
      end
      11'b10110111101 : begin
        result = input_1469;
      end
      11'b10110111110 : begin
        result = input_1470;
      end
      11'b10110111111 : begin
        result = input_1471;
      end
      11'b10111000000 : begin
        result = input_1472;
      end
      11'b10111000001 : begin
        result = input_1473;
      end
      11'b10111000010 : begin
        result = input_1474;
      end
      11'b10111000011 : begin
        result = input_1475;
      end
      11'b10111000100 : begin
        result = input_1476;
      end
      11'b10111000101 : begin
        result = input_1477;
      end
      11'b10111000110 : begin
        result = input_1478;
      end
      11'b10111000111 : begin
        result = input_1479;
      end
      11'b10111001000 : begin
        result = input_1480;
      end
      11'b10111001001 : begin
        result = input_1481;
      end
      11'b10111001010 : begin
        result = input_1482;
      end
      11'b10111001011 : begin
        result = input_1483;
      end
      11'b10111001100 : begin
        result = input_1484;
      end
      11'b10111001101 : begin
        result = input_1485;
      end
      11'b10111001110 : begin
        result = input_1486;
      end
      11'b10111001111 : begin
        result = input_1487;
      end
      11'b10111010000 : begin
        result = input_1488;
      end
      11'b10111010001 : begin
        result = input_1489;
      end
      11'b10111010010 : begin
        result = input_1490;
      end
      11'b10111010011 : begin
        result = input_1491;
      end
      11'b10111010100 : begin
        result = input_1492;
      end
      11'b10111010101 : begin
        result = input_1493;
      end
      11'b10111010110 : begin
        result = input_1494;
      end
      11'b10111010111 : begin
        result = input_1495;
      end
      11'b10111011000 : begin
        result = input_1496;
      end
      11'b10111011001 : begin
        result = input_1497;
      end
      11'b10111011010 : begin
        result = input_1498;
      end
      11'b10111011011 : begin
        result = input_1499;
      end
      11'b10111011100 : begin
        result = input_1500;
      end
      11'b10111011101 : begin
        result = input_1501;
      end
      11'b10111011110 : begin
        result = input_1502;
      end
      11'b10111011111 : begin
        result = input_1503;
      end
      11'b10111100000 : begin
        result = input_1504;
      end
      11'b10111100001 : begin
        result = input_1505;
      end
      11'b10111100010 : begin
        result = input_1506;
      end
      11'b10111100011 : begin
        result = input_1507;
      end
      11'b10111100100 : begin
        result = input_1508;
      end
      11'b10111100101 : begin
        result = input_1509;
      end
      11'b10111100110 : begin
        result = input_1510;
      end
      11'b10111100111 : begin
        result = input_1511;
      end
      11'b10111101000 : begin
        result = input_1512;
      end
      11'b10111101001 : begin
        result = input_1513;
      end
      11'b10111101010 : begin
        result = input_1514;
      end
      11'b10111101011 : begin
        result = input_1515;
      end
      11'b10111101100 : begin
        result = input_1516;
      end
      11'b10111101101 : begin
        result = input_1517;
      end
      11'b10111101110 : begin
        result = input_1518;
      end
      11'b10111101111 : begin
        result = input_1519;
      end
      11'b10111110000 : begin
        result = input_1520;
      end
      11'b10111110001 : begin
        result = input_1521;
      end
      11'b10111110010 : begin
        result = input_1522;
      end
      11'b10111110011 : begin
        result = input_1523;
      end
      11'b10111110100 : begin
        result = input_1524;
      end
      11'b10111110101 : begin
        result = input_1525;
      end
      11'b10111110110 : begin
        result = input_1526;
      end
      11'b10111110111 : begin
        result = input_1527;
      end
      11'b10111111000 : begin
        result = input_1528;
      end
      11'b10111111001 : begin
        result = input_1529;
      end
      11'b10111111010 : begin
        result = input_1530;
      end
      11'b10111111011 : begin
        result = input_1531;
      end
      11'b10111111100 : begin
        result = input_1532;
      end
      11'b10111111101 : begin
        result = input_1533;
      end
      11'b10111111110 : begin
        result = input_1534;
      end
      11'b10111111111 : begin
        result = input_1535;
      end
      11'b11000000000 : begin
        result = input_1536;
      end
      11'b11000000001 : begin
        result = input_1537;
      end
      11'b11000000010 : begin
        result = input_1538;
      end
      11'b11000000011 : begin
        result = input_1539;
      end
      11'b11000000100 : begin
        result = input_1540;
      end
      11'b11000000101 : begin
        result = input_1541;
      end
      11'b11000000110 : begin
        result = input_1542;
      end
      11'b11000000111 : begin
        result = input_1543;
      end
      11'b11000001000 : begin
        result = input_1544;
      end
      11'b11000001001 : begin
        result = input_1545;
      end
      11'b11000001010 : begin
        result = input_1546;
      end
      11'b11000001011 : begin
        result = input_1547;
      end
      11'b11000001100 : begin
        result = input_1548;
      end
      11'b11000001101 : begin
        result = input_1549;
      end
      11'b11000001110 : begin
        result = input_1550;
      end
      11'b11000001111 : begin
        result = input_1551;
      end
      11'b11000010000 : begin
        result = input_1552;
      end
      11'b11000010001 : begin
        result = input_1553;
      end
      11'b11000010010 : begin
        result = input_1554;
      end
      11'b11000010011 : begin
        result = input_1555;
      end
      11'b11000010100 : begin
        result = input_1556;
      end
      11'b11000010101 : begin
        result = input_1557;
      end
      11'b11000010110 : begin
        result = input_1558;
      end
      11'b11000010111 : begin
        result = input_1559;
      end
      11'b11000011000 : begin
        result = input_1560;
      end
      11'b11000011001 : begin
        result = input_1561;
      end
      11'b11000011010 : begin
        result = input_1562;
      end
      11'b11000011011 : begin
        result = input_1563;
      end
      11'b11000011100 : begin
        result = input_1564;
      end
      11'b11000011101 : begin
        result = input_1565;
      end
      11'b11000011110 : begin
        result = input_1566;
      end
      11'b11000011111 : begin
        result = input_1567;
      end
      11'b11000100000 : begin
        result = input_1568;
      end
      11'b11000100001 : begin
        result = input_1569;
      end
      11'b11000100010 : begin
        result = input_1570;
      end
      11'b11000100011 : begin
        result = input_1571;
      end
      11'b11000100100 : begin
        result = input_1572;
      end
      11'b11000100101 : begin
        result = input_1573;
      end
      11'b11000100110 : begin
        result = input_1574;
      end
      11'b11000100111 : begin
        result = input_1575;
      end
      11'b11000101000 : begin
        result = input_1576;
      end
      11'b11000101001 : begin
        result = input_1577;
      end
      11'b11000101010 : begin
        result = input_1578;
      end
      11'b11000101011 : begin
        result = input_1579;
      end
      11'b11000101100 : begin
        result = input_1580;
      end
      11'b11000101101 : begin
        result = input_1581;
      end
      11'b11000101110 : begin
        result = input_1582;
      end
      11'b11000101111 : begin
        result = input_1583;
      end
      11'b11000110000 : begin
        result = input_1584;
      end
      11'b11000110001 : begin
        result = input_1585;
      end
      11'b11000110010 : begin
        result = input_1586;
      end
      11'b11000110011 : begin
        result = input_1587;
      end
      11'b11000110100 : begin
        result = input_1588;
      end
      11'b11000110101 : begin
        result = input_1589;
      end
      11'b11000110110 : begin
        result = input_1590;
      end
      11'b11000110111 : begin
        result = input_1591;
      end
      11'b11000111000 : begin
        result = input_1592;
      end
      11'b11000111001 : begin
        result = input_1593;
      end
      11'b11000111010 : begin
        result = input_1594;
      end
      11'b11000111011 : begin
        result = input_1595;
      end
      11'b11000111100 : begin
        result = input_1596;
      end
      11'b11000111101 : begin
        result = input_1597;
      end
      11'b11000111110 : begin
        result = input_1598;
      end
      11'b11000111111 : begin
        result = input_1599;
      end
      11'b11001000000 : begin
        result = input_1600;
      end
      11'b11001000001 : begin
        result = input_1601;
      end
      11'b11001000010 : begin
        result = input_1602;
      end
      11'b11001000011 : begin
        result = input_1603;
      end
      11'b11001000100 : begin
        result = input_1604;
      end
      11'b11001000101 : begin
        result = input_1605;
      end
      11'b11001000110 : begin
        result = input_1606;
      end
      11'b11001000111 : begin
        result = input_1607;
      end
      11'b11001001000 : begin
        result = input_1608;
      end
      11'b11001001001 : begin
        result = input_1609;
      end
      11'b11001001010 : begin
        result = input_1610;
      end
      11'b11001001011 : begin
        result = input_1611;
      end
      11'b11001001100 : begin
        result = input_1612;
      end
      11'b11001001101 : begin
        result = input_1613;
      end
      11'b11001001110 : begin
        result = input_1614;
      end
      11'b11001001111 : begin
        result = input_1615;
      end
      11'b11001010000 : begin
        result = input_1616;
      end
      11'b11001010001 : begin
        result = input_1617;
      end
      11'b11001010010 : begin
        result = input_1618;
      end
      11'b11001010011 : begin
        result = input_1619;
      end
      11'b11001010100 : begin
        result = input_1620;
      end
      11'b11001010101 : begin
        result = input_1621;
      end
      11'b11001010110 : begin
        result = input_1622;
      end
      11'b11001010111 : begin
        result = input_1623;
      end
      11'b11001011000 : begin
        result = input_1624;
      end
      11'b11001011001 : begin
        result = input_1625;
      end
      11'b11001011010 : begin
        result = input_1626;
      end
      11'b11001011011 : begin
        result = input_1627;
      end
      11'b11001011100 : begin
        result = input_1628;
      end
      11'b11001011101 : begin
        result = input_1629;
      end
      11'b11001011110 : begin
        result = input_1630;
      end
      11'b11001011111 : begin
        result = input_1631;
      end
      11'b11001100000 : begin
        result = input_1632;
      end
      11'b11001100001 : begin
        result = input_1633;
      end
      11'b11001100010 : begin
        result = input_1634;
      end
      11'b11001100011 : begin
        result = input_1635;
      end
      11'b11001100100 : begin
        result = input_1636;
      end
      11'b11001100101 : begin
        result = input_1637;
      end
      11'b11001100110 : begin
        result = input_1638;
      end
      11'b11001100111 : begin
        result = input_1639;
      end
      11'b11001101000 : begin
        result = input_1640;
      end
      11'b11001101001 : begin
        result = input_1641;
      end
      11'b11001101010 : begin
        result = input_1642;
      end
      11'b11001101011 : begin
        result = input_1643;
      end
      11'b11001101100 : begin
        result = input_1644;
      end
      11'b11001101101 : begin
        result = input_1645;
      end
      11'b11001101110 : begin
        result = input_1646;
      end
      11'b11001101111 : begin
        result = input_1647;
      end
      11'b11001110000 : begin
        result = input_1648;
      end
      11'b11001110001 : begin
        result = input_1649;
      end
      11'b11001110010 : begin
        result = input_1650;
      end
      11'b11001110011 : begin
        result = input_1651;
      end
      11'b11001110100 : begin
        result = input_1652;
      end
      11'b11001110101 : begin
        result = input_1653;
      end
      11'b11001110110 : begin
        result = input_1654;
      end
      11'b11001110111 : begin
        result = input_1655;
      end
      11'b11001111000 : begin
        result = input_1656;
      end
      11'b11001111001 : begin
        result = input_1657;
      end
      11'b11001111010 : begin
        result = input_1658;
      end
      11'b11001111011 : begin
        result = input_1659;
      end
      11'b11001111100 : begin
        result = input_1660;
      end
      11'b11001111101 : begin
        result = input_1661;
      end
      11'b11001111110 : begin
        result = input_1662;
      end
      11'b11001111111 : begin
        result = input_1663;
      end
      11'b11010000000 : begin
        result = input_1664;
      end
      11'b11010000001 : begin
        result = input_1665;
      end
      11'b11010000010 : begin
        result = input_1666;
      end
      11'b11010000011 : begin
        result = input_1667;
      end
      11'b11010000100 : begin
        result = input_1668;
      end
      11'b11010000101 : begin
        result = input_1669;
      end
      11'b11010000110 : begin
        result = input_1670;
      end
      11'b11010000111 : begin
        result = input_1671;
      end
      11'b11010001000 : begin
        result = input_1672;
      end
      11'b11010001001 : begin
        result = input_1673;
      end
      11'b11010001010 : begin
        result = input_1674;
      end
      11'b11010001011 : begin
        result = input_1675;
      end
      11'b11010001100 : begin
        result = input_1676;
      end
      11'b11010001101 : begin
        result = input_1677;
      end
      11'b11010001110 : begin
        result = input_1678;
      end
      11'b11010001111 : begin
        result = input_1679;
      end
      11'b11010010000 : begin
        result = input_1680;
      end
      11'b11010010001 : begin
        result = input_1681;
      end
      11'b11010010010 : begin
        result = input_1682;
      end
      11'b11010010011 : begin
        result = input_1683;
      end
      11'b11010010100 : begin
        result = input_1684;
      end
      11'b11010010101 : begin
        result = input_1685;
      end
      11'b11010010110 : begin
        result = input_1686;
      end
      11'b11010010111 : begin
        result = input_1687;
      end
      11'b11010011000 : begin
        result = input_1688;
      end
      11'b11010011001 : begin
        result = input_1689;
      end
      11'b11010011010 : begin
        result = input_1690;
      end
      11'b11010011011 : begin
        result = input_1691;
      end
      11'b11010011100 : begin
        result = input_1692;
      end
      11'b11010011101 : begin
        result = input_1693;
      end
      11'b11010011110 : begin
        result = input_1694;
      end
      11'b11010011111 : begin
        result = input_1695;
      end
      11'b11010100000 : begin
        result = input_1696;
      end
      11'b11010100001 : begin
        result = input_1697;
      end
      11'b11010100010 : begin
        result = input_1698;
      end
      11'b11010100011 : begin
        result = input_1699;
      end
      11'b11010100100 : begin
        result = input_1700;
      end
      11'b11010100101 : begin
        result = input_1701;
      end
      11'b11010100110 : begin
        result = input_1702;
      end
      11'b11010100111 : begin
        result = input_1703;
      end
      11'b11010101000 : begin
        result = input_1704;
      end
      11'b11010101001 : begin
        result = input_1705;
      end
      11'b11010101010 : begin
        result = input_1706;
      end
      11'b11010101011 : begin
        result = input_1707;
      end
      11'b11010101100 : begin
        result = input_1708;
      end
      11'b11010101101 : begin
        result = input_1709;
      end
      11'b11010101110 : begin
        result = input_1710;
      end
      11'b11010101111 : begin
        result = input_1711;
      end
      11'b11010110000 : begin
        result = input_1712;
      end
      11'b11010110001 : begin
        result = input_1713;
      end
      11'b11010110010 : begin
        result = input_1714;
      end
      11'b11010110011 : begin
        result = input_1715;
      end
      11'b11010110100 : begin
        result = input_1716;
      end
      11'b11010110101 : begin
        result = input_1717;
      end
      11'b11010110110 : begin
        result = input_1718;
      end
      11'b11010110111 : begin
        result = input_1719;
      end
      11'b11010111000 : begin
        result = input_1720;
      end
      11'b11010111001 : begin
        result = input_1721;
      end
      11'b11010111010 : begin
        result = input_1722;
      end
      11'b11010111011 : begin
        result = input_1723;
      end
      11'b11010111100 : begin
        result = input_1724;
      end
      11'b11010111101 : begin
        result = input_1725;
      end
      11'b11010111110 : begin
        result = input_1726;
      end
      11'b11010111111 : begin
        result = input_1727;
      end
      11'b11011000000 : begin
        result = input_1728;
      end
      11'b11011000001 : begin
        result = input_1729;
      end
      11'b11011000010 : begin
        result = input_1730;
      end
      11'b11011000011 : begin
        result = input_1731;
      end
      11'b11011000100 : begin
        result = input_1732;
      end
      11'b11011000101 : begin
        result = input_1733;
      end
      11'b11011000110 : begin
        result = input_1734;
      end
      11'b11011000111 : begin
        result = input_1735;
      end
      11'b11011001000 : begin
        result = input_1736;
      end
      11'b11011001001 : begin
        result = input_1737;
      end
      11'b11011001010 : begin
        result = input_1738;
      end
      11'b11011001011 : begin
        result = input_1739;
      end
      11'b11011001100 : begin
        result = input_1740;
      end
      11'b11011001101 : begin
        result = input_1741;
      end
      11'b11011001110 : begin
        result = input_1742;
      end
      11'b11011001111 : begin
        result = input_1743;
      end
      11'b11011010000 : begin
        result = input_1744;
      end
      11'b11011010001 : begin
        result = input_1745;
      end
      11'b11011010010 : begin
        result = input_1746;
      end
      11'b11011010011 : begin
        result = input_1747;
      end
      11'b11011010100 : begin
        result = input_1748;
      end
      11'b11011010101 : begin
        result = input_1749;
      end
      11'b11011010110 : begin
        result = input_1750;
      end
      11'b11011010111 : begin
        result = input_1751;
      end
      11'b11011011000 : begin
        result = input_1752;
      end
      11'b11011011001 : begin
        result = input_1753;
      end
      11'b11011011010 : begin
        result = input_1754;
      end
      11'b11011011011 : begin
        result = input_1755;
      end
      11'b11011011100 : begin
        result = input_1756;
      end
      11'b11011011101 : begin
        result = input_1757;
      end
      11'b11011011110 : begin
        result = input_1758;
      end
      11'b11011011111 : begin
        result = input_1759;
      end
      11'b11011100000 : begin
        result = input_1760;
      end
      11'b11011100001 : begin
        result = input_1761;
      end
      11'b11011100010 : begin
        result = input_1762;
      end
      11'b11011100011 : begin
        result = input_1763;
      end
      11'b11011100100 : begin
        result = input_1764;
      end
      11'b11011100101 : begin
        result = input_1765;
      end
      11'b11011100110 : begin
        result = input_1766;
      end
      11'b11011100111 : begin
        result = input_1767;
      end
      11'b11011101000 : begin
        result = input_1768;
      end
      11'b11011101001 : begin
        result = input_1769;
      end
      11'b11011101010 : begin
        result = input_1770;
      end
      11'b11011101011 : begin
        result = input_1771;
      end
      11'b11011101100 : begin
        result = input_1772;
      end
      11'b11011101101 : begin
        result = input_1773;
      end
      11'b11011101110 : begin
        result = input_1774;
      end
      11'b11011101111 : begin
        result = input_1775;
      end
      11'b11011110000 : begin
        result = input_1776;
      end
      11'b11011110001 : begin
        result = input_1777;
      end
      11'b11011110010 : begin
        result = input_1778;
      end
      11'b11011110011 : begin
        result = input_1779;
      end
      11'b11011110100 : begin
        result = input_1780;
      end
      11'b11011110101 : begin
        result = input_1781;
      end
      11'b11011110110 : begin
        result = input_1782;
      end
      11'b11011110111 : begin
        result = input_1783;
      end
      11'b11011111000 : begin
        result = input_1784;
      end
      11'b11011111001 : begin
        result = input_1785;
      end
      11'b11011111010 : begin
        result = input_1786;
      end
      11'b11011111011 : begin
        result = input_1787;
      end
      11'b11011111100 : begin
        result = input_1788;
      end
      11'b11011111101 : begin
        result = input_1789;
      end
      11'b11011111110 : begin
        result = input_1790;
      end
      default : begin
        result = input_1791;
      end
    endcase
    MUX_v_5_1792_2 = result;
  end
  endfunction

endmodule




//------> ./myproject_ROM_1i9_1o5_e071483337062336669c4105b16859e3bb.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
//
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Mon Oct 24 20:35:20 2022
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i9_1o5_e071483337062336669c4105b16859e3bb
// ------------------------------------------------------------------


module converterBlock_ROM_1i9_1o5_e071483337062336669c4105b16859e3bb (
  I_1, O_1
);
  input [8:0] I_1;
  output [4:0] O_1;



  // Interconnect Declarations for Component Instantiations
  assign O_1 = MUX_v_5_384_2(5'b11111, 5'b10111, 5'b01010, 5'b11111, 5'b10101, 5'b01010,
      5'b11010, 5'b01011, 5'b10000, 5'b11111, 5'b01111, 5'b10000, 5'b00011, 5'b10101,
      5'b01100, 5'b11100, 5'b11100, 5'b00100, 5'b11111, 5'b11110, 5'b01010, 5'b00100,
      5'b01000, 5'b10101, 5'b11100, 5'b10111, 5'b01110, 5'b00100, 5'b01001, 5'b10000,
      5'b00010, 5'b11001, 5'b00111, 5'b11101, 5'b01010, 5'b10010, 5'b00000, 5'b11011,
      5'b11110, 5'b11011, 5'b01001, 5'b11001, 5'b11110, 5'b01100, 5'b10110, 5'b00010,
      5'b11000, 5'b00100, 5'b00110, 5'b10111, 5'b00000, 5'b00011, 5'b11111, 5'b11110,
      5'b11000, 5'b00110, 5'b11100, 5'b00100, 5'b10110, 5'b01010, 5'b11111, 5'b01011,
      5'b10011, 5'b11101, 5'b00110, 5'b10101, 5'b00001, 5'b10111, 5'b01010, 5'b00000,
      5'b10100, 5'b01001, 5'b11011, 5'b01010, 5'b11001, 5'b11101, 5'b01100, 5'b10110,
      5'b00010, 5'b10111, 5'b00010, 5'b00001, 5'b01101, 5'b10000, 5'b00001, 5'b01010,
      5'b10111, 5'b11111, 5'b01110, 5'b10000, 5'b00000, 5'b11001, 5'b01000, 5'b00001,
      5'b11100, 5'b01001, 5'b11101, 5'b00011, 5'b00011, 5'b00101, 5'b10100, 5'b01000,
      5'b11101, 5'b00011, 5'b00110, 5'b00101, 5'b00000, 5'b11011, 5'b00011, 5'b11011,
      5'b00011, 5'b00011, 5'b00011, 5'b10111, 5'b11001, 5'b11111, 5'b01010, 5'b01001,
      5'b00000, 5'b10101, 5'b00011, 5'b11101, 5'b11101, 5'b00100, 5'b00101, 5'b10110,
      5'b11101, 5'b11011, 5'b01000, 5'b11101, 5'b01111, 5'b10000, 5'b11011, 5'b11000,
      5'b01001, 5'b10111, 5'b00100, 5'b00000, 5'b11100, 5'b01100, 5'b10110, 5'b11111,
      5'b01100, 5'b10100, 5'b00011, 5'b00100, 5'b11000, 5'b11110, 5'b11001, 5'b00100,
      5'b11110, 5'b01001, 5'b10111, 5'b00001, 5'b01100, 5'b11000, 5'b11111, 5'b10101,
      5'b00101, 5'b11111, 5'b01110, 5'b10010, 5'b11111, 5'b10111, 5'b01000, 5'b11110,
      5'b11010, 5'b01010, 5'b00010, 5'b01100, 5'b10001, 5'b00100, 5'b00110, 5'b11000,
      5'b00001, 5'b01100, 5'b10000, 5'b00001, 5'b01011, 5'b10110, 5'b00010, 5'b10011,
      5'b01010, 5'b00001, 5'b10010, 5'b01010, 5'b00100, 5'b00111, 5'b11010, 5'b11100,
      5'b11111, 5'b01000, 5'b11111, 5'b01111, 5'b10000, 5'b11001, 5'b01011, 5'b10111,
      5'b10110, 5'b00010, 5'b00001, 5'b11011, 5'b11000, 5'b01011, 5'b00010, 5'b11001,
      5'b01000, 5'b00101, 5'b11101, 5'b11010, 5'b00010, 5'b10111, 5'b01010, 5'b11111,
      5'b01101, 5'b10100, 5'b00010, 5'b01100, 5'b10101, 5'b00001, 5'b01001, 5'b10101,
      5'b00100, 5'b01010, 5'b10111, 5'b11110, 5'b01100, 5'b10000, 5'b11101, 5'b11101,
      5'b01000, 5'b11111, 5'b01100, 5'b10011, 5'b11111, 5'b11100, 5'b00111, 5'b11110,
      5'b11110, 5'b00100, 5'b00000, 5'b11011, 5'b00110, 5'b00010, 5'b01010, 5'b10110,
      5'b11111, 5'b00110, 5'b10000, 5'b00100, 5'b00110, 5'b10101, 5'b00011, 5'b01011,
      5'b10000, 5'b00001, 5'b10110, 5'b01011, 5'b01001, 5'b11011, 5'b00010, 5'b11001,
      5'b10101, 5'b01100, 5'b11010, 5'b11100, 5'b00100, 5'b11111, 5'b00110, 5'b10111,
      5'b00000, 5'b00111, 5'b10101, 5'b00010, 5'b10001, 5'b00111, 5'b11110, 5'b01111,
      5'b10001, 5'b00000, 5'b11000, 5'b01001, 5'b11100, 5'b11110, 5'b00101, 5'b11101,
      5'b00110, 5'b11011, 5'b11011, 5'b00100, 5'b00001, 5'b11011, 5'b01001, 5'b11001,
      5'b11100, 5'b01010, 5'b10000, 5'b00001, 5'b11001, 5'b01010, 5'b00010, 5'b01001,
      5'b10100, 5'b11110, 5'b01100, 5'b10000, 5'b11100, 5'b01111, 5'b10001, 5'b00000,
      5'b11101, 5'b00111, 5'b00000, 5'b10101, 5'b01100, 5'b11101, 5'b10011, 5'b01000,
      5'b11100, 5'b11111, 5'b00100, 5'b11111, 5'b01000, 5'b11001, 5'b11111, 5'b01000,
      5'b11011, 5'b10111, 5'b00110, 5'b11011, 5'b00011, 5'b11101, 5'b11111, 5'b11111,
      5'b01011, 5'b10101, 5'b00100, 5'b11010, 5'b00101, 5'b00110, 5'b10100, 5'b00110,
      5'b00010, 5'b00110, 5'b11001, 5'b11100, 5'b00011, 5'b00011, 5'b00010, 5'b01000,
      5'b10011, 5'b01001, 5'b11101, 5'b11101, 5'b11110, 5'b01011, 5'b10000, 5'b11010,
      5'b01010, 5'b11001, 5'b00110, 5'b00010, 5'b11000, 5'b01001, 5'b10110, 5'b01010,
      5'b11101, 5'b01111, 5'b10000, 5'b00100, 5'b10111, 5'b01011, 5'b00001, 5'b01011,
      5'b10100, 5'b11110, 5'b01011, 5'b10101, 5'b00000, 5'b01000, 5'b10101, 5'b11111,
      5'b11010, 5'b01101, I_1);

  function automatic [4:0] MUX_v_5_384_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [4:0] input_4;
    input [4:0] input_5;
    input [4:0] input_6;
    input [4:0] input_7;
    input [4:0] input_8;
    input [4:0] input_9;
    input [4:0] input_10;
    input [4:0] input_11;
    input [4:0] input_12;
    input [4:0] input_13;
    input [4:0] input_14;
    input [4:0] input_15;
    input [4:0] input_16;
    input [4:0] input_17;
    input [4:0] input_18;
    input [4:0] input_19;
    input [4:0] input_20;
    input [4:0] input_21;
    input [4:0] input_22;
    input [4:0] input_23;
    input [4:0] input_24;
    input [4:0] input_25;
    input [4:0] input_26;
    input [4:0] input_27;
    input [4:0] input_28;
    input [4:0] input_29;
    input [4:0] input_30;
    input [4:0] input_31;
    input [4:0] input_32;
    input [4:0] input_33;
    input [4:0] input_34;
    input [4:0] input_35;
    input [4:0] input_36;
    input [4:0] input_37;
    input [4:0] input_38;
    input [4:0] input_39;
    input [4:0] input_40;
    input [4:0] input_41;
    input [4:0] input_42;
    input [4:0] input_43;
    input [4:0] input_44;
    input [4:0] input_45;
    input [4:0] input_46;
    input [4:0] input_47;
    input [4:0] input_48;
    input [4:0] input_49;
    input [4:0] input_50;
    input [4:0] input_51;
    input [4:0] input_52;
    input [4:0] input_53;
    input [4:0] input_54;
    input [4:0] input_55;
    input [4:0] input_56;
    input [4:0] input_57;
    input [4:0] input_58;
    input [4:0] input_59;
    input [4:0] input_60;
    input [4:0] input_61;
    input [4:0] input_62;
    input [4:0] input_63;
    input [4:0] input_64;
    input [4:0] input_65;
    input [4:0] input_66;
    input [4:0] input_67;
    input [4:0] input_68;
    input [4:0] input_69;
    input [4:0] input_70;
    input [4:0] input_71;
    input [4:0] input_72;
    input [4:0] input_73;
    input [4:0] input_74;
    input [4:0] input_75;
    input [4:0] input_76;
    input [4:0] input_77;
    input [4:0] input_78;
    input [4:0] input_79;
    input [4:0] input_80;
    input [4:0] input_81;
    input [4:0] input_82;
    input [4:0] input_83;
    input [4:0] input_84;
    input [4:0] input_85;
    input [4:0] input_86;
    input [4:0] input_87;
    input [4:0] input_88;
    input [4:0] input_89;
    input [4:0] input_90;
    input [4:0] input_91;
    input [4:0] input_92;
    input [4:0] input_93;
    input [4:0] input_94;
    input [4:0] input_95;
    input [4:0] input_96;
    input [4:0] input_97;
    input [4:0] input_98;
    input [4:0] input_99;
    input [4:0] input_100;
    input [4:0] input_101;
    input [4:0] input_102;
    input [4:0] input_103;
    input [4:0] input_104;
    input [4:0] input_105;
    input [4:0] input_106;
    input [4:0] input_107;
    input [4:0] input_108;
    input [4:0] input_109;
    input [4:0] input_110;
    input [4:0] input_111;
    input [4:0] input_112;
    input [4:0] input_113;
    input [4:0] input_114;
    input [4:0] input_115;
    input [4:0] input_116;
    input [4:0] input_117;
    input [4:0] input_118;
    input [4:0] input_119;
    input [4:0] input_120;
    input [4:0] input_121;
    input [4:0] input_122;
    input [4:0] input_123;
    input [4:0] input_124;
    input [4:0] input_125;
    input [4:0] input_126;
    input [4:0] input_127;
    input [4:0] input_128;
    input [4:0] input_129;
    input [4:0] input_130;
    input [4:0] input_131;
    input [4:0] input_132;
    input [4:0] input_133;
    input [4:0] input_134;
    input [4:0] input_135;
    input [4:0] input_136;
    input [4:0] input_137;
    input [4:0] input_138;
    input [4:0] input_139;
    input [4:0] input_140;
    input [4:0] input_141;
    input [4:0] input_142;
    input [4:0] input_143;
    input [4:0] input_144;
    input [4:0] input_145;
    input [4:0] input_146;
    input [4:0] input_147;
    input [4:0] input_148;
    input [4:0] input_149;
    input [4:0] input_150;
    input [4:0] input_151;
    input [4:0] input_152;
    input [4:0] input_153;
    input [4:0] input_154;
    input [4:0] input_155;
    input [4:0] input_156;
    input [4:0] input_157;
    input [4:0] input_158;
    input [4:0] input_159;
    input [4:0] input_160;
    input [4:0] input_161;
    input [4:0] input_162;
    input [4:0] input_163;
    input [4:0] input_164;
    input [4:0] input_165;
    input [4:0] input_166;
    input [4:0] input_167;
    input [4:0] input_168;
    input [4:0] input_169;
    input [4:0] input_170;
    input [4:0] input_171;
    input [4:0] input_172;
    input [4:0] input_173;
    input [4:0] input_174;
    input [4:0] input_175;
    input [4:0] input_176;
    input [4:0] input_177;
    input [4:0] input_178;
    input [4:0] input_179;
    input [4:0] input_180;
    input [4:0] input_181;
    input [4:0] input_182;
    input [4:0] input_183;
    input [4:0] input_184;
    input [4:0] input_185;
    input [4:0] input_186;
    input [4:0] input_187;
    input [4:0] input_188;
    input [4:0] input_189;
    input [4:0] input_190;
    input [4:0] input_191;
    input [4:0] input_192;
    input [4:0] input_193;
    input [4:0] input_194;
    input [4:0] input_195;
    input [4:0] input_196;
    input [4:0] input_197;
    input [4:0] input_198;
    input [4:0] input_199;
    input [4:0] input_200;
    input [4:0] input_201;
    input [4:0] input_202;
    input [4:0] input_203;
    input [4:0] input_204;
    input [4:0] input_205;
    input [4:0] input_206;
    input [4:0] input_207;
    input [4:0] input_208;
    input [4:0] input_209;
    input [4:0] input_210;
    input [4:0] input_211;
    input [4:0] input_212;
    input [4:0] input_213;
    input [4:0] input_214;
    input [4:0] input_215;
    input [4:0] input_216;
    input [4:0] input_217;
    input [4:0] input_218;
    input [4:0] input_219;
    input [4:0] input_220;
    input [4:0] input_221;
    input [4:0] input_222;
    input [4:0] input_223;
    input [4:0] input_224;
    input [4:0] input_225;
    input [4:0] input_226;
    input [4:0] input_227;
    input [4:0] input_228;
    input [4:0] input_229;
    input [4:0] input_230;
    input [4:0] input_231;
    input [4:0] input_232;
    input [4:0] input_233;
    input [4:0] input_234;
    input [4:0] input_235;
    input [4:0] input_236;
    input [4:0] input_237;
    input [4:0] input_238;
    input [4:0] input_239;
    input [4:0] input_240;
    input [4:0] input_241;
    input [4:0] input_242;
    input [4:0] input_243;
    input [4:0] input_244;
    input [4:0] input_245;
    input [4:0] input_246;
    input [4:0] input_247;
    input [4:0] input_248;
    input [4:0] input_249;
    input [4:0] input_250;
    input [4:0] input_251;
    input [4:0] input_252;
    input [4:0] input_253;
    input [4:0] input_254;
    input [4:0] input_255;
    input [4:0] input_256;
    input [4:0] input_257;
    input [4:0] input_258;
    input [4:0] input_259;
    input [4:0] input_260;
    input [4:0] input_261;
    input [4:0] input_262;
    input [4:0] input_263;
    input [4:0] input_264;
    input [4:0] input_265;
    input [4:0] input_266;
    input [4:0] input_267;
    input [4:0] input_268;
    input [4:0] input_269;
    input [4:0] input_270;
    input [4:0] input_271;
    input [4:0] input_272;
    input [4:0] input_273;
    input [4:0] input_274;
    input [4:0] input_275;
    input [4:0] input_276;
    input [4:0] input_277;
    input [4:0] input_278;
    input [4:0] input_279;
    input [4:0] input_280;
    input [4:0] input_281;
    input [4:0] input_282;
    input [4:0] input_283;
    input [4:0] input_284;
    input [4:0] input_285;
    input [4:0] input_286;
    input [4:0] input_287;
    input [4:0] input_288;
    input [4:0] input_289;
    input [4:0] input_290;
    input [4:0] input_291;
    input [4:0] input_292;
    input [4:0] input_293;
    input [4:0] input_294;
    input [4:0] input_295;
    input [4:0] input_296;
    input [4:0] input_297;
    input [4:0] input_298;
    input [4:0] input_299;
    input [4:0] input_300;
    input [4:0] input_301;
    input [4:0] input_302;
    input [4:0] input_303;
    input [4:0] input_304;
    input [4:0] input_305;
    input [4:0] input_306;
    input [4:0] input_307;
    input [4:0] input_308;
    input [4:0] input_309;
    input [4:0] input_310;
    input [4:0] input_311;
    input [4:0] input_312;
    input [4:0] input_313;
    input [4:0] input_314;
    input [4:0] input_315;
    input [4:0] input_316;
    input [4:0] input_317;
    input [4:0] input_318;
    input [4:0] input_319;
    input [4:0] input_320;
    input [4:0] input_321;
    input [4:0] input_322;
    input [4:0] input_323;
    input [4:0] input_324;
    input [4:0] input_325;
    input [4:0] input_326;
    input [4:0] input_327;
    input [4:0] input_328;
    input [4:0] input_329;
    input [4:0] input_330;
    input [4:0] input_331;
    input [4:0] input_332;
    input [4:0] input_333;
    input [4:0] input_334;
    input [4:0] input_335;
    input [4:0] input_336;
    input [4:0] input_337;
    input [4:0] input_338;
    input [4:0] input_339;
    input [4:0] input_340;
    input [4:0] input_341;
    input [4:0] input_342;
    input [4:0] input_343;
    input [4:0] input_344;
    input [4:0] input_345;
    input [4:0] input_346;
    input [4:0] input_347;
    input [4:0] input_348;
    input [4:0] input_349;
    input [4:0] input_350;
    input [4:0] input_351;
    input [4:0] input_352;
    input [4:0] input_353;
    input [4:0] input_354;
    input [4:0] input_355;
    input [4:0] input_356;
    input [4:0] input_357;
    input [4:0] input_358;
    input [4:0] input_359;
    input [4:0] input_360;
    input [4:0] input_361;
    input [4:0] input_362;
    input [4:0] input_363;
    input [4:0] input_364;
    input [4:0] input_365;
    input [4:0] input_366;
    input [4:0] input_367;
    input [4:0] input_368;
    input [4:0] input_369;
    input [4:0] input_370;
    input [4:0] input_371;
    input [4:0] input_372;
    input [4:0] input_373;
    input [4:0] input_374;
    input [4:0] input_375;
    input [4:0] input_376;
    input [4:0] input_377;
    input [4:0] input_378;
    input [4:0] input_379;
    input [4:0] input_380;
    input [4:0] input_381;
    input [4:0] input_382;
    input [4:0] input_383;
    input [8:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      9'b101000011 : begin
        result = input_323;
      end
      9'b101000100 : begin
        result = input_324;
      end
      9'b101000101 : begin
        result = input_325;
      end
      9'b101000110 : begin
        result = input_326;
      end
      9'b101000111 : begin
        result = input_327;
      end
      9'b101001000 : begin
        result = input_328;
      end
      9'b101001001 : begin
        result = input_329;
      end
      9'b101001010 : begin
        result = input_330;
      end
      9'b101001011 : begin
        result = input_331;
      end
      9'b101001100 : begin
        result = input_332;
      end
      9'b101001101 : begin
        result = input_333;
      end
      9'b101001110 : begin
        result = input_334;
      end
      9'b101001111 : begin
        result = input_335;
      end
      9'b101010000 : begin
        result = input_336;
      end
      9'b101010001 : begin
        result = input_337;
      end
      9'b101010010 : begin
        result = input_338;
      end
      9'b101010011 : begin
        result = input_339;
      end
      9'b101010100 : begin
        result = input_340;
      end
      9'b101010101 : begin
        result = input_341;
      end
      9'b101010110 : begin
        result = input_342;
      end
      9'b101010111 : begin
        result = input_343;
      end
      9'b101011000 : begin
        result = input_344;
      end
      9'b101011001 : begin
        result = input_345;
      end
      9'b101011010 : begin
        result = input_346;
      end
      9'b101011011 : begin
        result = input_347;
      end
      9'b101011100 : begin
        result = input_348;
      end
      9'b101011101 : begin
        result = input_349;
      end
      9'b101011110 : begin
        result = input_350;
      end
      9'b101011111 : begin
        result = input_351;
      end
      9'b101100000 : begin
        result = input_352;
      end
      9'b101100001 : begin
        result = input_353;
      end
      9'b101100010 : begin
        result = input_354;
      end
      9'b101100011 : begin
        result = input_355;
      end
      9'b101100100 : begin
        result = input_356;
      end
      9'b101100101 : begin
        result = input_357;
      end
      9'b101100110 : begin
        result = input_358;
      end
      9'b101100111 : begin
        result = input_359;
      end
      9'b101101000 : begin
        result = input_360;
      end
      9'b101101001 : begin
        result = input_361;
      end
      9'b101101010 : begin
        result = input_362;
      end
      9'b101101011 : begin
        result = input_363;
      end
      9'b101101100 : begin
        result = input_364;
      end
      9'b101101101 : begin
        result = input_365;
      end
      9'b101101110 : begin
        result = input_366;
      end
      9'b101101111 : begin
        result = input_367;
      end
      9'b101110000 : begin
        result = input_368;
      end
      9'b101110001 : begin
        result = input_369;
      end
      9'b101110010 : begin
        result = input_370;
      end
      9'b101110011 : begin
        result = input_371;
      end
      9'b101110100 : begin
        result = input_372;
      end
      9'b101110101 : begin
        result = input_373;
      end
      9'b101110110 : begin
        result = input_374;
      end
      9'b101110111 : begin
        result = input_375;
      end
      9'b101111000 : begin
        result = input_376;
      end
      9'b101111001 : begin
        result = input_377;
      end
      9'b101111010 : begin
        result = input_378;
      end
      9'b101111011 : begin
        result = input_379;
      end
      9'b101111100 : begin
        result = input_380;
      end
      9'b101111101 : begin
        result = input_381;
      end
      9'b101111110 : begin
        result = input_382;
      end
      default : begin
        result = input_383;
      end
    endcase
    MUX_v_5_384_2 = result;
  end
  endfunction

endmodule




//------> ./myproject.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
// 
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Mon Oct 24 20:58:28 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module converterBlock_myproject_core_core_fsm (
  clk, rst, fsm_output, Product2_C_0_tr0, Product1_C_1_tr0, Accum2_C_0_tr0, Accum1_C_0_tr0,
      Product2_1_C_0_tr0, Result_C_3_tr0, Accum2_1_C_0_tr0, Accum1_1_C_0_tr0, Result_1_C_1_tr0
);
  input clk;
  input rst;
  output [14:0] fsm_output;
  reg [14:0] fsm_output;
  input Product2_C_0_tr0;
  input Product1_C_1_tr0;
  input Accum2_C_0_tr0;
  input Accum1_C_0_tr0;
  input Product2_1_C_0_tr0;
  input Result_C_3_tr0;
  input Accum2_1_C_0_tr0;
  input Accum1_1_C_0_tr0;
  input Result_1_C_1_tr0;


  // FSM State Type Declaration for converterBlock_myproject_core_core_fsm_1
  parameter
    main_C_0 = 4'd0,
    Product1_C_0 = 4'd1,
    Product2_C_0 = 4'd2,
    Product1_C_1 = 4'd3,
    Accum2_C_0 = 4'd4,
    Accum1_C_0 = 4'd5,
    Result_C_0 = 4'd6,
    Result_C_1 = 4'd7,
    Result_C_2 = 4'd8,
    Product2_1_C_0 = 4'd9,
    Result_C_3 = 4'd10,
    Accum2_1_C_0 = 4'd11,
    Accum1_1_C_0 = 4'd12,
    Result_1_C_0 = 4'd13,
    Result_1_C_1 = 4'd14;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : converterBlock_myproject_core_core_fsm_1
    case (state_var)
      Product1_C_0 : begin
        fsm_output = 15'b000000000000010;
        state_var_NS = Product2_C_0;
      end
      Product2_C_0 : begin
        fsm_output = 15'b000000000000100;
        if ( Product2_C_0_tr0 ) begin
          state_var_NS = Product1_C_1;
        end
        else begin
          state_var_NS = Product2_C_0;
        end
      end
      Product1_C_1 : begin
        fsm_output = 15'b000000000001000;
        if ( Product1_C_1_tr0 ) begin
          state_var_NS = Accum2_C_0;
        end
        else begin
          state_var_NS = Product1_C_0;
        end
      end
      Accum2_C_0 : begin
        fsm_output = 15'b000000000010000;
        if ( Accum2_C_0_tr0 ) begin
          state_var_NS = Accum1_C_0;
        end
        else begin
          state_var_NS = Accum2_C_0;
        end
      end
      Accum1_C_0 : begin
        fsm_output = 15'b000000000100000;
        if ( Accum1_C_0_tr0 ) begin
          state_var_NS = Result_C_0;
        end
        else begin
          state_var_NS = Accum2_C_0;
        end
      end
      Result_C_0 : begin
        fsm_output = 15'b000000001000000;
        state_var_NS = Result_C_1;
      end
      Result_C_1 : begin
        fsm_output = 15'b000000010000000;
        state_var_NS = Result_C_2;
      end
      Result_C_2 : begin
        fsm_output = 15'b000000100000000;
        state_var_NS = Product2_1_C_0;
      end
      Product2_1_C_0 : begin
        fsm_output = 15'b000001000000000;
        if ( Product2_1_C_0_tr0 ) begin
          state_var_NS = Result_C_3;
        end
        else begin
          state_var_NS = Product2_1_C_0;
        end
      end
      Result_C_3 : begin
        fsm_output = 15'b000010000000000;
        if ( Result_C_3_tr0 ) begin
          state_var_NS = Accum2_1_C_0;
        end
        else begin
          state_var_NS = Result_C_0;
        end
      end
      Accum2_1_C_0 : begin
        fsm_output = 15'b000100000000000;
        if ( Accum2_1_C_0_tr0 ) begin
          state_var_NS = Accum1_1_C_0;
        end
        else begin
          state_var_NS = Accum2_1_C_0;
        end
      end
      Accum1_1_C_0 : begin
        fsm_output = 15'b001000000000000;
        if ( Accum1_1_C_0_tr0 ) begin
          state_var_NS = Result_1_C_0;
        end
        else begin
          state_var_NS = Accum2_1_C_0;
        end
      end
      Result_1_C_0 : begin
        fsm_output = 15'b010000000000000;
        state_var_NS = Result_1_C_1;
      end
      Result_1_C_1 : begin
        fsm_output = 15'b100000000000000;
        if ( Result_1_C_1_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = Result_1_C_0;
        end
      end
      // main_C_0
      default : begin
        fsm_output = 15'b000000000000001;
        state_var_NS = Product1_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core
// ------------------------------------------------------------------


module converterBlock_myproject_core (
  clk, rst, input_1_rsc_dat, layer6_out_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer6_out_rsc_dat;


  // Interconnect Declarations
  wire [223:0] input_1_rsci_idat;
  reg [15:0] layer6_out_rsci_idat_47_32;
  reg [15:0] layer6_out_rsci_idat_31_16;
  reg [15:0] layer6_out_rsci_idat_15_0;
  wire [14:0] fsm_output;
  wire Result_and_1_tmp;
  wire or_dcpl_69;
  wire or_dcpl_70;
  wire or_dcpl_80;
  wire or_dcpl_81;
  wire or_dcpl_420;
  wire or_dcpl_423;
  wire or_dcpl_682;
  wire or_dcpl_683;
  wire or_dcpl_686;
  wire or_dcpl_687;
  wire or_dcpl_946;
  wire or_dcpl_949;
  wire and_dcpl_2;
  wire or_dcpl_2015;
  wire or_dcpl_2016;
  wire or_dcpl_2020;
  wire or_dcpl_2027;
  wire or_dcpl_2028;
  wire or_dcpl_2029;
  wire or_dcpl_2030;
  wire or_dcpl_2031;
  wire or_dcpl_2032;
  wire or_dcpl_2035;
  wire or_dcpl_2037;
  wire or_dcpl_2038;
  wire or_dcpl_2040;
  wire or_dcpl_2041;
  wire or_dcpl_2042;
  wire or_dcpl_2043;
  wire or_dcpl_2045;
  wire or_dcpl_2046;
  wire or_dcpl_2047;
  wire or_dcpl_2048;
  wire or_dcpl_2049;
  wire or_dcpl_2050;
  wire or_dcpl_2052;
  wire or_dcpl_2053;
  wire or_dcpl_2054;
  wire or_dcpl_2057;
  wire or_dcpl_2059;
  wire or_dcpl_2060;
  wire or_dcpl_2062;
  wire or_dcpl_2063;
  wire or_dcpl_2064;
  wire or_dcpl_2066;
  wire or_dcpl_2067;
  wire or_dcpl_2069;
  wire or_dcpl_2070;
  wire or_dcpl_2072;
  wire or_dcpl_2074;
  wire or_dcpl_2076;
  wire or_dcpl_2078;
  wire or_dcpl_2079;
  wire or_dcpl_2080;
  wire or_dcpl_2081;
  wire or_dcpl_2083;
  wire or_dcpl_2085;
  wire or_dcpl_2087;
  wire or_dcpl_2089;
  wire or_dcpl_2093;
  wire or_dcpl_2095;
  wire or_dcpl_2107;
  wire or_dcpl_2110;
  wire or_dcpl_2112;
  wire or_dcpl_2113;
  wire or_dcpl_2115;
  wire or_dcpl_2117;
  wire or_dcpl_2120;
  wire or_dcpl_2122;
  wire or_dcpl_2124;
  wire or_dcpl_2126;
  wire or_dcpl_2129;
  wire or_dcpl_2131;
  wire or_dcpl_2133;
  wire or_dcpl_2135;
  wire or_dcpl_2137;
  wire or_dcpl_2140;
  wire or_dcpl_2141;
  wire or_dcpl_2142;
  wire or_dcpl_2160;
  wire or_dcpl_2179;
  wire or_dcpl_2180;
  wire or_dcpl_2234;
  wire or_dcpl_2273;
  wire or_dcpl_2291;
  wire or_dcpl_2310;
  wire or_dcpl_2330;
  wire or_dcpl_2419;
  wire or_dcpl_2423;
  wire or_dcpl_2441;
  wire or_dcpl_2461;
  wire or_dcpl_2479;
  wire or_dcpl_2570;
  wire or_dcpl_2589;
  wire or_dcpl_2607;
  wire or_dcpl_2609;
  wire or_dcpl_2627;
  wire or_dcpl_2717;
  wire or_dcpl_2718;
  wire or_dcpl_2737;
  wire or_dcpl_2738;
  wire or_dcpl_2756;
  wire or_dcpl_2775;
  wire or_dcpl_2793;
  wire or_dcpl_2795;
  wire or_dcpl_2867;
  wire or_dcpl_2886;
  wire or_dcpl_2904;
  wire or_dcpl_2924;
  wire or_dcpl_2977;
  wire or_dcpl_3100;
  wire or_dcpl_3119;
  wire or_dcpl_3137;
  wire or_dcpl_3157;
  wire or_dcpl_3246;
  wire or_dcpl_3266;
  wire or_dcpl_3284;
  wire or_dcpl_3303;
  wire or_dcpl_3393;
  wire or_dcpl_3411;
  wire or_dcpl_3430;
  wire or_dcpl_3449;
  wire or_dcpl_3539;
  wire or_dcpl_3557;
  wire or_dcpl_3576;
  wire or_dcpl_3594;
  wire or_dcpl_3684;
  wire or_dcpl_3703;
  wire or_dcpl_3723;
  wire or_dcpl_3741;
  wire or_dcpl_3830;
  wire or_dcpl_3850;
  wire or_dcpl_3947;
  wire or_dcpl_3948;
  wire or_dcpl_3949;
  wire or_dcpl_3950;
  wire or_dcpl_3951;
  wire or_dcpl_3952;
  wire or_dcpl_3953;
  wire or_dcpl_3955;
  wire or_dcpl_3956;
  wire or_dcpl_3958;
  wire or_dcpl_3959;
  wire or_dcpl_3960;
  wire or_dcpl_3962;
  wire or_dcpl_3963;
  wire or_dcpl_3964;
  wire or_dcpl_3965;
  wire or_dcpl_3966;
  wire or_dcpl_3968;
  wire or_dcpl_3969;
  wire or_dcpl_3971;
  wire or_dcpl_3974;
  wire or_dcpl_3979;
  wire or_dcpl_3980;
  wire or_dcpl_3984;
  wire or_dcpl_3987;
  wire or_dcpl_3988;
  wire or_dcpl_3990;
  wire or_dcpl_3992;
  wire or_dcpl_4008;
  wire or_dcpl_4009;
  wire or_dcpl_4010;
  wire or_dcpl_4014;
  wire or_dcpl_4015;
  wire or_dcpl_4018;
  wire or_dcpl_4021;
  wire or_dcpl_4024;
  wire or_dcpl_4027;
  wire or_dcpl_4031;
  wire or_dcpl_4034;
  wire or_dcpl_4037;
  wire or_dcpl_4038;
  wire or_dcpl_4040;
  wire or_dcpl_4058;
  wire or_dcpl_4060;
  wire or_dcpl_4077;
  wire or_dcpl_4079;
  wire or_dcpl_4097;
  wire or_dcpl_4099;
  wire or_dcpl_4117;
  wire or_dcpl_4119;
  wire or_dcpl_4172;
  wire or_dcpl_4173;
  wire or_dcpl_4174;
  wire or_dcpl_4177;
  wire or_dcpl_4178;
  wire or_dcpl_4182;
  wire or_dcpl_4185;
  wire or_dcpl_4188;
  wire or_dcpl_4191;
  wire or_dcpl_4194;
  wire or_dcpl_4198;
  wire or_dcpl_4396;
  wire or_dcpl_4397;
  wire or_dcpl_4398;
  wire or_dcpl_4399;
  wire and_dcpl_20;
  wire and_dcpl_21;
  wire and_dcpl_22;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire or_dcpl_4409;
  wire or_dcpl_4410;
  wire or_dcpl_4411;
  wire or_dcpl_4412;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire or_dcpl_4414;
  wire or_dcpl_4415;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire or_dcpl_4419;
  wire or_dcpl_4420;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire or_dcpl_4422;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire or_dcpl_4424;
  wire and_dcpl_56;
  wire or_dcpl_4428;
  wire and_dcpl_58;
  wire or_dcpl_4430;
  wire and_dcpl_60;
  wire or_dcpl_4432;
  wire and_dcpl_62;
  wire or_dcpl_4434;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire or_dcpl_4456;
  wire or_dcpl_4457;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire or_dcpl_4459;
  wire or_dcpl_4460;
  wire and_dcpl_93;
  wire or_dcpl_4464;
  wire and_dcpl_95;
  wire or_dcpl_4466;
  wire and_dcpl_123;
  wire or_dcpl_4494;
  wire and_dcpl_125;
  wire or_dcpl_4496;
  wire and_dcpl_129;
  wire or_dcpl_4500;
  wire and_dcpl_131;
  wire or_dcpl_4502;
  wire and_dcpl_159;
  wire or_dcpl_4530;
  wire and_dcpl_161;
  wire or_dcpl_4532;
  wire and_dcpl_165;
  wire or_dcpl_4536;
  wire and_dcpl_167;
  wire or_dcpl_4538;
  wire or_tmp_2362;
  wire or_tmp_2754;
  wire and_5035_cse;
  wire and_5068_cse;
  reg Result_1_Result_1_nor_itm;
  wire [15:0] Accum2_mux_131;
  reg [3:0] Accum1_ii_3_0_sva;
  reg [7:0] nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1;
  reg [7:0] Result_ires_7_0_sva_1;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_0_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_1_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_2_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_3_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_4_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_5_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_6_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_7_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_8_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_9_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_10_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_11_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_12_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_13_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_14_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_15_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_16_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_17_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_18_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_19_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_20_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_21_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_22_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_23_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_24_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_25_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_26_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_27_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_28_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_29_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_30_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_31_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_32_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_33_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_34_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_35_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_36_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_37_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_38_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_39_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_40_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_41_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_42_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_43_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_44_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_45_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_46_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_47_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_48_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_49_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_50_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_51_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_52_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_53_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_54_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_55_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_56_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_57_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_58_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_59_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_60_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_61_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_62_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_63_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_64_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_65_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_66_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_67_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_68_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_69_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_70_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_71_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_72_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_73_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_74_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_75_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_76_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_77_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_78_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_79_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_80_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_81_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_82_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_83_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_84_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_85_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_86_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_87_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_88_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_89_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_90_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_91_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_92_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_93_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_94_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_95_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_96_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_97_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_98_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_99_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_100_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_101_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_102_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_103_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_104_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_105_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_106_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_107_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_108_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_109_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_110_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_111_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_112_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_113_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_114_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_115_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_116_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_117_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_118_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_119_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_120_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_121_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_122_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_123_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_124_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_125_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_126_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_127_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_128_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_129_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_130_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_131_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_132_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_133_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_134_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_135_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_136_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_137_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_138_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_139_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_140_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_141_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_142_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_143_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_144_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_145_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_146_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_147_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_148_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_149_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_150_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_151_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_152_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_153_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_154_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_155_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_156_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_157_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_158_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_159_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_160_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_161_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_162_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_163_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_164_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_165_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_166_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_167_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_168_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_169_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_170_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_171_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_172_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_173_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_174_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_175_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_176_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_177_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_178_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_179_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_180_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_181_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_182_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_183_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_184_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_185_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_186_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_187_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_188_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_189_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_190_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_191_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_192_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_193_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_194_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_195_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_196_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_197_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_198_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_199_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_200_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_201_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_202_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_203_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_204_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_205_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_206_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_207_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_208_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_209_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_210_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_211_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_212_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_213_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_214_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_215_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_216_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_217_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_218_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_219_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_220_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_221_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_222_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_223_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_224_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_225_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_226_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_227_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_228_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_229_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_230_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_231_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_232_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_233_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_234_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_235_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_236_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_237_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_238_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_239_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_240_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_241_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_242_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_243_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_244_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_245_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_246_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_247_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_248_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_249_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_250_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_251_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_252_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_253_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_254_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_255_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_256_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_257_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_258_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_259_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_260_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_261_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_262_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_263_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_264_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_265_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_266_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_267_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_268_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_269_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_270_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_271_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_272_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_273_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_274_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_275_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_276_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_277_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_278_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_279_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_280_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_281_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_282_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_283_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_284_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_285_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_286_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_287_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_288_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_289_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_290_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_291_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_292_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_293_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_294_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_295_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_296_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_297_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_298_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_299_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_300_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_301_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_302_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_303_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_304_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_305_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_306_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_307_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_308_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_309_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_310_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_311_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_312_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_313_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_314_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_315_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_316_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_317_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_318_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_319_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_320_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_321_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_322_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_323_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_324_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_325_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_326_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_327_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_328_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_329_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_330_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_331_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_332_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_333_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_334_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_335_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_336_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_337_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_338_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_339_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_340_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_341_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_342_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_343_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_344_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_345_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_346_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_347_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_348_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_349_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_350_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_351_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_352_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_353_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_354_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_355_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_356_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_357_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_358_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_359_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_360_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_361_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_362_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_363_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_364_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_365_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_366_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_367_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_368_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_369_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_370_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_371_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_372_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_373_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_374_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_375_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_376_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_377_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_378_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_379_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_380_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_381_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_382_reg;
  reg [10:0] reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_383_reg;
  wire [3:0] z_out;
  wire [4:0] nl_z_out;
  wire [3:0] z_out_1;
  wire [4:0] nl_z_out_1;
  wire [7:0] z_out_2;
  wire [8:0] nl_z_out_2;
  wire [15:0] z_out_6;
  wire [16:0] nl_z_out_6;
  reg [15:0] nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_31_16_lpi_2;
  reg [15:0] nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_47_32_lpi_2;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_895_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_896_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_894_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_897_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_893_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_898_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_892_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_899_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_891_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_900_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_890_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_901_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_889_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_902_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_888_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_903_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_887_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_904_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_886_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_905_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_885_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_906_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_884_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_907_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_883_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_908_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_882_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_909_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_881_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_910_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_880_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_911_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_879_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_912_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_878_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_913_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_877_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_914_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_876_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_915_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_875_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_916_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_874_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_917_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_873_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_918_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_872_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_919_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_871_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_920_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_870_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_921_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_869_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_922_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_868_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_923_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_867_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_924_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_866_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_925_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_865_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_926_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_864_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_927_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_863_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_928_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_862_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_929_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_861_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_930_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_860_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_931_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_859_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_932_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_858_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_933_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_857_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_934_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_856_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_935_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_855_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_936_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_854_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_937_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_853_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_938_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_852_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_939_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_851_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_940_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_850_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_941_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_849_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_942_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_848_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_943_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_847_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_944_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_846_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_945_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_845_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_946_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_844_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_947_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_843_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_948_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_842_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_949_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_841_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_950_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_840_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_951_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_839_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_952_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_838_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_953_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_837_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_954_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_836_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_955_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_835_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_956_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_834_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_957_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_833_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_958_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_832_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_959_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_831_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_960_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_830_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_961_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_829_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_962_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_828_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_963_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_827_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_964_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_826_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_965_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_825_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_966_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_824_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_967_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_823_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_968_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_822_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_969_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_821_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_970_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_820_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_971_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_819_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_972_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_818_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_973_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_817_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_974_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_816_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_975_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_815_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_976_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_814_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_977_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_813_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_978_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_812_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_979_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_811_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_980_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_810_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_981_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_809_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_982_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_808_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_983_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_807_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_984_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_806_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_985_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_805_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_986_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_804_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_987_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_803_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_988_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_802_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_989_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_801_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_990_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_800_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_991_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_799_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_992_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_798_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_993_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_797_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_994_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_796_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_995_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_795_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_996_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_794_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_997_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_793_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_998_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_792_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_999_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_791_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1000_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_790_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1001_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_789_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1002_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_788_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1003_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_787_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1004_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_786_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1005_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_785_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1006_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_784_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1007_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_783_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1008_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_782_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1009_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_781_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1010_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_780_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1011_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_779_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1012_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_778_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1013_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_777_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1014_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_776_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1015_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_775_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1016_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_774_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1017_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_773_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1018_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_772_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1019_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_771_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1020_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_770_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1021_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_769_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1022_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_768_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1023_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_767_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1024_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_766_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1025_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_765_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1026_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_764_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1027_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_763_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1028_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_762_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1029_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_761_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1030_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_760_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1031_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_759_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1032_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_758_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1033_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_757_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1034_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_756_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1035_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_755_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1036_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_754_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1037_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_753_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1038_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_752_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1039_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_751_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1040_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_750_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1041_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_749_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1042_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_748_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1043_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_747_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1044_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_746_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1045_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_745_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1046_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_744_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1047_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_743_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1048_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_742_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1049_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_741_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1050_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_740_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1051_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_739_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1052_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_738_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1053_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_737_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1054_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_736_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1055_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_735_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1056_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_734_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1057_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_733_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1058_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_732_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1059_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_731_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1060_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_730_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1061_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_729_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1062_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_728_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1063_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_727_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1064_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_726_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1065_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_725_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1066_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_724_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1067_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_723_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1068_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_722_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1069_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_721_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1070_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_720_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1071_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_719_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1072_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_718_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1073_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_717_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1074_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_716_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1075_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_715_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1076_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_714_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1077_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_713_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1078_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_712_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1079_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_711_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1080_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_710_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1081_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_709_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1082_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_708_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1083_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_707_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1084_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_706_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1085_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_705_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1086_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_704_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1087_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_703_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1088_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_702_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1089_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_701_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1090_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_700_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1091_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_699_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1092_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_698_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1093_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_697_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1094_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_696_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1095_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_695_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1096_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_694_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1097_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_693_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1098_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_692_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1099_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_691_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1100_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_690_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1101_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_689_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1102_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_688_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1103_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_687_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1104_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_686_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1105_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_685_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1106_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_684_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1107_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_683_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1108_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_682_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1109_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_681_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1110_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_680_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1111_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_679_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1112_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_678_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1113_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_677_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1114_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_676_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1115_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_675_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1116_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_674_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1117_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_673_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1118_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_672_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1119_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_671_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1120_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_670_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1121_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_669_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1122_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_668_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1123_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_667_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1124_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_666_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1125_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_665_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1126_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_664_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1127_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_663_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1128_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_662_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1129_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_661_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1130_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_660_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1131_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_659_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1132_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_658_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1133_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_657_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1134_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_656_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1135_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_655_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1136_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_654_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1137_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_653_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1138_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_652_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1139_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_651_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1140_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_650_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1141_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_649_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1142_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_648_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1143_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_647_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1144_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_646_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1145_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_645_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1146_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_644_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1147_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_643_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1148_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_642_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1149_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_641_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1150_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_640_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1151_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_639_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1152_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_638_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1153_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_637_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1154_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_636_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1155_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_635_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1156_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_634_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1157_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_633_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1158_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_632_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1159_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_631_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1160_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_630_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1161_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_629_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1162_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_628_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1163_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_627_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1164_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_626_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1165_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_625_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1166_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_624_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1167_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_623_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1168_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_622_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1169_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_621_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1170_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_620_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1171_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_619_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1172_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_618_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1173_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_617_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1174_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_616_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1175_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_615_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1176_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_614_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1177_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_613_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1178_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_612_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1179_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_611_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1180_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_610_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1181_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_609_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1182_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_608_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1183_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_607_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1184_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_606_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1185_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_605_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1186_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_604_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1187_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_603_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1188_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_602_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1189_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_601_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1190_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_600_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1191_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_599_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1192_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_598_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1193_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_597_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1194_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_596_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1195_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_595_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1196_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_594_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1197_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_593_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1198_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_592_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1199_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_591_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1200_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_590_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1201_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_589_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1202_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_588_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1203_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_587_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1204_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_586_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1205_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_585_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1206_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_584_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1207_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_583_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1208_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_582_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1209_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_581_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1210_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_580_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1211_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_579_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1212_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_578_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1213_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_577_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1214_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_576_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1215_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_575_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1216_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_574_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1217_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_573_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1218_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_572_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1219_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_571_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1220_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_570_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1221_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_569_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1222_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_568_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1223_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_567_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1224_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_566_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1225_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_565_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1226_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_564_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1227_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_563_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1228_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_562_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1229_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_561_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1230_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_560_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1231_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_559_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1232_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_558_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1233_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_557_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1234_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_556_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1235_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_555_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1236_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_554_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1237_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_553_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1238_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_552_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1239_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_551_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1240_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_550_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1241_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_549_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1242_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_548_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1243_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_547_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1244_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_546_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1245_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_545_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1246_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_544_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1247_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_543_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1248_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_542_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1249_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_541_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1250_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_540_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1251_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_539_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1252_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_538_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1253_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_537_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1254_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_536_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1255_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_535_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1256_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_534_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1257_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_533_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1258_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_532_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1259_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_531_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1260_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_530_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1261_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_529_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1262_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_528_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1263_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_527_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1264_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_526_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1265_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_525_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1266_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_524_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1267_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_523_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1268_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_522_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1269_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_521_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1270_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_520_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1271_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_519_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1272_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_518_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1273_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_517_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1274_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_516_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1275_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_515_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1276_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_514_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1277_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_513_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1278_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_512_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1279_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_511_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1280_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_510_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1281_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_509_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1282_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_508_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1283_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_507_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1284_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_506_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1285_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_505_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1286_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_504_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1287_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_503_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1288_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_502_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1289_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_501_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1290_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_500_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1291_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_499_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1292_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_498_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1293_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_497_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1294_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_496_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1295_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_495_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1296_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_494_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1297_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_493_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1298_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_492_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1299_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_491_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1300_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_490_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1301_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_489_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1302_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_488_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1303_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_487_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1304_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_486_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1305_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_485_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1306_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_484_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1307_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_483_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1308_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_482_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1309_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_481_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1310_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_480_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1311_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_479_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1312_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_478_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1313_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_477_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1314_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_476_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1315_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_475_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1316_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_474_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1317_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_473_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1318_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_472_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1319_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_471_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1320_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_470_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1321_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_469_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1322_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_468_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1323_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_467_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1324_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_466_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1325_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_465_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1326_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_464_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1327_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_463_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1328_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_462_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1329_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_461_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1330_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_460_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1331_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_459_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1332_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_458_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1333_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_457_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1334_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_456_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1335_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_455_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1336_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_454_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1337_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_453_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1338_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_452_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1339_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_451_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1340_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_450_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1341_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_449_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1342_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_448_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1343_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_447_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1344_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_446_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1345_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_445_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1346_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_444_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1347_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_443_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1348_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_442_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1349_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_441_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1350_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_440_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1351_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_439_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1352_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_438_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1353_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_437_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1354_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_436_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1355_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_435_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1356_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_434_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1357_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_433_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1358_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_432_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1359_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_431_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1360_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_430_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1361_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_429_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1362_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_428_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1363_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_427_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1364_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_426_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1365_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_425_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1366_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_424_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1367_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_423_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1368_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_422_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1369_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_421_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1370_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_420_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1371_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_419_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1372_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_418_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1373_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_417_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1374_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_416_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1375_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_415_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1376_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_414_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1377_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_413_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1378_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_412_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1379_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_411_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1380_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_410_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1381_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_409_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1382_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_408_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1383_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_407_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1384_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_406_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1385_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_405_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1386_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_404_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1387_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_403_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1388_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_402_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1389_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_401_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1390_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_400_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1391_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_399_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1392_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_398_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1393_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_397_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1394_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_396_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1395_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_395_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1396_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_394_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1397_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_393_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1398_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_392_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1399_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_391_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1400_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_390_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1401_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_389_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1402_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_388_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1403_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_387_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1404_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_386_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1405_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_385_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1406_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_384_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1407_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_383_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1408_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_382_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1409_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_381_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1410_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_380_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1411_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_379_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1412_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_378_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1413_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_377_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1414_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_376_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1415_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_375_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1416_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_374_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1417_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_373_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1418_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_372_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1419_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_371_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1420_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_370_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1421_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_369_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1422_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_368_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1423_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_367_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1424_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_366_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1425_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_365_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1426_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_364_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1427_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_363_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1428_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_362_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1429_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_361_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1430_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_360_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1431_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_359_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1432_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_358_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1433_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_357_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1434_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_356_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1435_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_355_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1436_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_354_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1437_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_353_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1438_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_352_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1439_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_351_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1440_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_350_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1441_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_349_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1442_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_348_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1443_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_347_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1444_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_346_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1445_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_345_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1446_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_344_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1447_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_343_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1448_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_342_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1449_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_341_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1450_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_340_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1451_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_339_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1452_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_338_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1453_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_337_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1454_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_336_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1455_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_335_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1456_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_334_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1457_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_333_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1458_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_332_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1459_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_331_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1460_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_330_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1461_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_329_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1462_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_328_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1463_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_327_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1464_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_326_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1465_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_325_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1466_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_324_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1467_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_323_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1468_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_322_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1469_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_321_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1470_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_320_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1471_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_319_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1472_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_318_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1473_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_317_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1474_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_316_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1475_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_315_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1476_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_314_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1477_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_313_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1478_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_312_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1479_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_311_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1480_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_310_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1481_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_309_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1482_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_308_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1483_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_307_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1484_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_306_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1485_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_305_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1486_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_304_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1487_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_303_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1488_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_302_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1489_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_301_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1490_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_300_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1491_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_299_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1492_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_298_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1493_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_297_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1494_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_296_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1495_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_295_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1496_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_294_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1497_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_293_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1498_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_292_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1499_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_291_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1500_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_290_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1501_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_289_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1502_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_288_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1503_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_287_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1504_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_286_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1505_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_285_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1506_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_284_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1507_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_283_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1508_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_282_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1509_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_281_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1510_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_280_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1511_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_279_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1512_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_278_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1513_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_277_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1514_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_276_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1515_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_275_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1516_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_274_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1517_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_273_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1518_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_272_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1519_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_271_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1520_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_270_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1521_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_269_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1522_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_268_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1523_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_267_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1524_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_266_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1525_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_265_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1526_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_264_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1527_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_263_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1528_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_262_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1529_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_261_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1530_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_260_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1531_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_259_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1532_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_258_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1533_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_257_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1534_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_256_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1535_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_255_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1536_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_254_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1537_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_253_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1538_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_252_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1539_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_251_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1540_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_250_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1541_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_249_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1542_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_248_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1543_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_247_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1544_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_246_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1545_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_245_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1546_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_244_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1547_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_243_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1548_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_242_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1549_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_241_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1550_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_240_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1551_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_239_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1552_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_238_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1553_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_237_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1554_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_236_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1555_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_235_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1556_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_234_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1557_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_233_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1558_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_232_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1559_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_231_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1560_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_230_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1561_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_229_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1562_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_228_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1563_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_227_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1564_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_226_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1565_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_225_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1566_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_224_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1567_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_223_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1568_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_222_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1569_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_221_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1570_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_220_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1571_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_219_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1572_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_218_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1573_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_217_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1574_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_216_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1575_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_215_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1576_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_214_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1577_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_213_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1578_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_212_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1579_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_211_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1580_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_210_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1581_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_209_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1582_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_208_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1583_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_207_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1584_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_206_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1585_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_205_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1586_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_204_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1587_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_203_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1588_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_202_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1589_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_201_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1590_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_200_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1591_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_199_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1592_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_198_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1593_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_197_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1594_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_196_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1595_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_195_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1596_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_194_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1597_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_193_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1598_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_192_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1599_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_191_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1600_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_190_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1601_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_189_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1602_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_188_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1603_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_187_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1604_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_186_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1605_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_185_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1606_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_184_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1607_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_183_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1608_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_182_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1609_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_181_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1610_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_180_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1611_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_179_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1612_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_178_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1613_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_177_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1614_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_176_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1615_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_175_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1616_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_174_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1617_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_173_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1618_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_172_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1619_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_171_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1620_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_170_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1621_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_169_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1622_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_168_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1623_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_167_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1624_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_166_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1625_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_165_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1626_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_164_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1627_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_163_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1628_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_162_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1629_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_161_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1630_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_160_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1631_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_159_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1632_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_158_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1633_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_157_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1634_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_156_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1635_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_155_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1636_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_154_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1637_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_153_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1638_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_152_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1639_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_151_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1640_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_150_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1641_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_149_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1642_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_148_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1643_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_147_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1644_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_146_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1645_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_145_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1646_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_144_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1647_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_143_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1648_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_142_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1649_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_141_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1650_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_140_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1651_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_139_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1652_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_138_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1653_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_137_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1654_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_136_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1655_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_135_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1656_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_134_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1657_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_133_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1658_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_132_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1659_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_131_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1660_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_130_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1661_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_129_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1662_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_128_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1663_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_127_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1664_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_126_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1665_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_125_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1666_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_124_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1667_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_123_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1668_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_122_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1669_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_121_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1670_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_120_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1671_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_119_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1672_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_118_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1673_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_117_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1674_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_116_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1675_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_115_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1676_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_114_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1677_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_113_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1678_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_112_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1679_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_111_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1680_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_110_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1681_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_109_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1682_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_108_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1683_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_107_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1684_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_106_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1685_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_105_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1686_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_104_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1687_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_103_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1688_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_102_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1689_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_101_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1690_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_100_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1691_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_99_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1692_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_98_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1693_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_97_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1694_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_96_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1695_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_95_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1696_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_94_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1697_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_93_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1698_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_92_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1699_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_91_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1700_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_90_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1701_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_89_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1702_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_88_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1703_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_87_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1704_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_86_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1705_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_85_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1706_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_84_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1707_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_83_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1708_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_82_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1709_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_81_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1710_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_80_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1711_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_79_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1712_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_78_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1713_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_77_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1714_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_76_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1715_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_75_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1716_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_74_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1717_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_73_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1718_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_72_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1719_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_71_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1720_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_70_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1721_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_69_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1722_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_68_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1723_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_67_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1724_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_66_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1725_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_65_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1726_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_64_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1727_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_63_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1728_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_62_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1729_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_61_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1730_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_60_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1731_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_59_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1732_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_58_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1733_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_57_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1734_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_56_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1735_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_55_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1736_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_54_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1737_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_53_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1738_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_52_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1739_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_51_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1740_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_50_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1741_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_49_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1742_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_48_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1743_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_47_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1744_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_46_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1745_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_45_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1746_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_44_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1747_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_43_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1748_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_42_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1749_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_41_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1750_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_40_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1751_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_39_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1752_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_38_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1753_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_37_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1754_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_36_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1755_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_35_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1756_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_34_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1757_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_33_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1758_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_32_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1759_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_31_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1760_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_30_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1761_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_29_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1762_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_28_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1763_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_27_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1764_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_26_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1765_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_25_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1766_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_24_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1767_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_23_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1768_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_22_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1769_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_21_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1770_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_20_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1771_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_19_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1772_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_18_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1773_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_17_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1774_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_16_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1775_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_15_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1776_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_14_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1777_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_13_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1778_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_12_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1779_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_11_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1780_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_10_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1781_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_9_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1782_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_8_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1783_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_7_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1784_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_6_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1785_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_5_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1786_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_4_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1787_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_3_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1788_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_2_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1789_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1790_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_0_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_mult_1791_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_63_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_64_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_62_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_65_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_61_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_66_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_60_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_67_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_59_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_68_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_58_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_69_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_57_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_70_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_56_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_71_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_55_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_72_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_54_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_73_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_53_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_74_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_52_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_75_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_51_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_76_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_50_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_77_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_49_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_78_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_48_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_79_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_47_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_80_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_46_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_81_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_45_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_82_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_44_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_83_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_43_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_84_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_42_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_85_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_41_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_86_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_40_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_87_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_39_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_88_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_38_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_89_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_37_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_90_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_36_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_91_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_35_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_92_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_34_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_93_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_33_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_94_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_32_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_95_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_31_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_96_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_30_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_97_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_29_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_98_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_28_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_99_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_27_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_100_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_26_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_101_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_25_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_102_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_24_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_103_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_23_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_104_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_22_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_105_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_21_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_106_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_20_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_107_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_19_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_108_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_18_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_109_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_17_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_110_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_16_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_111_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_15_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_112_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_14_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_113_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_13_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_114_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_12_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_115_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_11_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_116_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_10_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_117_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_9_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_118_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_8_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_119_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_7_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_120_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_6_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_121_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_5_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_122_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_4_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_123_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_3_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_124_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_2_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_125_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_1_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_126_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_0_lpi_3;
  reg [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_127_lpi_3;
  reg layer4_out_9_lpi_2_dfm;
  reg [7:0] layer4_out_8_1_lpi_2_dfm;
  reg layer4_out_0_lpi_2_dfm;
  reg [7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_7_0_sva_1;
  reg [6:0] Product1_1_ii_7_0_sva_6_0;
  wire Accum1_ii_3_0_sva_mx0c0;
  wire Accum1_ii_3_0_sva_mx0c3;
  wire nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1_mx0c2;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1;
  wire [15:0] Accum2_1_mux_6;
  wire [4:0] ROM_1i11_1o5_815f6a3dbd0daa2d77beb65dd6cecbbc31_1;
  wire [4:0] ROM_1i9_1o5_4a143e9cb1f27bd26e0331874cec74ad2f_1;
  wire and_5052_rgt;
  wire or_6921_rgt;
  wire and_5057_rgt;
  wire and_5081_rgt;
  wire and_5086_rgt;
  wire and_5214_rgt;
  wire and_5219_rgt;
  wire Product1_1_ii_or_cse;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_or_cse;
  wire [15:0] nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
  wire [6:0] Product2_1_index_mux_cse;
  wire or_7342_cse;
  wire operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
  wire [15:0] z_out_5_19_4;
  wire [7:0] Product2_1_index_acc_sdt;
  wire [8:0] nl_Product2_1_index_acc_sdt;
  wire [7:0] z_out_4_8_1;
  wire [8:0] nl_z_out_4_8_1;

  wire and_655_nl;
  wire and_661_nl;
  wire and_667_nl;
  wire[3:0] Product1_ii_Product1_ii_mux_nl;
  wire[1:0] Product2_1_jj_Product2_1_jj_and_nl;
  wire[1:0] Product2_1_jj_mux_nl;
  wire nand_22_nl;
  wire Accum1_ii_not_1_nl;
  wire[15:0] Product1_mux_nl;
  wire nnet_dense_latency_input_t_layer2_t_config2_acc_or_nl;
  wire[6:0] mux_nl;
  wire[6:0] Product2_jj_and_nl;
  wire nor_23_nl;
  wire or_7339_nl;
  wire and_5067_nl;
  wire and_5074_nl;
  wire nnet_dense_latency_input_t_layer2_t_config2_acc_or_4_nl;
  wire and_5095_nl;
  wire and_5102_nl;
  wire and_5109_nl;
  wire and_5116_nl;
  wire and_5123_nl;
  wire and_5130_nl;
  wire and_5137_nl;
  wire and_5144_nl;
  wire and_5151_nl;
  wire and_5158_nl;
  wire and_5165_nl;
  wire and_5172_nl;
  wire and_5179_nl;
  wire and_5186_nl;
  wire and_5193_nl;
  wire and_5200_nl;
  wire and_5207_nl;
  wire nnet_dense_latency_input_t_layer2_t_config2_acc_or_23_nl;
  wire and_5228_nl;
  wire and_5235_nl;
  wire and_5242_nl;
  wire and_5249_nl;
  wire and_5256_nl;
  wire and_5263_nl;
  wire and_5270_nl;
  wire and_5277_nl;
  wire and_5284_nl;
  wire and_5291_nl;
  wire and_5298_nl;
  wire and_5305_nl;
  wire not_2388_nl;
  wire and_5319_nl;
  wire and_5333_nl;
  wire and_5340_nl;
  wire and_5354_nl;
  wire and_5361_nl;
  wire and_5368_nl;
  wire and_5375_nl;
  wire and_5382_nl;
  wire and_5389_nl;
  wire and_5396_nl;
  wire and_5403_nl;
  wire and_5410_nl;
  wire and_5417_nl;
  wire and_5424_nl;
  wire and_5431_nl;
  wire and_5438_nl;
  wire and_5445_nl;
  wire and_5452_nl;
  wire and_5461_nl;
  wire and_5468_nl;
  wire and_5475_nl;
  wire and_5482_nl;
  wire and_5489_nl;
  wire and_5496_nl;
  wire and_5503_nl;
  wire and_5510_nl;
  wire and_5517_nl;
  wire and_5524_nl;
  wire and_5531_nl;
  wire and_5538_nl;
  wire and_5545_nl;
  wire and_5552_nl;
  wire and_5559_nl;
  wire and_5566_nl;
  wire and_5580_nl;
  wire and_5587_nl;
  wire and_5594_nl;
  wire and_5601_nl;
  wire and_5608_nl;
  wire and_5615_nl;
  wire and_5629_nl;
  wire and_5636_nl;
  wire and_5643_nl;
  wire and_5650_nl;
  wire and_5657_nl;
  wire and_5664_nl;
  wire and_5671_nl;
  wire and_5678_nl;
  wire and_5685_nl;
  wire and_5692_nl;
  wire and_5699_nl;
  wire and_5706_nl;
  wire and_5713_nl;
  wire and_5720_nl;
  wire and_5727_nl;
  wire and_5734_nl;
  wire and_5741_nl;
  wire and_5748_nl;
  wire and_5755_nl;
  wire and_5769_nl;
  wire and_5776_nl;
  wire and_5783_nl;
  wire and_5790_nl;
  wire and_5797_nl;
  wire and_5804_nl;
  wire and_5811_nl;
  wire and_5818_nl;
  wire and_5825_nl;
  wire and_5832_nl;
  wire and_5839_nl;
  wire and_5846_nl;
  wire and_5853_nl;
  wire and_5860_nl;
  wire and_5867_nl;
  wire and_5874_nl;
  wire and_5881_nl;
  wire and_5888_nl;
  wire and_5895_nl;
  wire and_5902_nl;
  wire and_5909_nl;
  wire and_5916_nl;
  wire and_5923_nl;
  wire and_5930_nl;
  wire and_5937_nl;
  wire and_5944_nl;
  wire and_5951_nl;
  wire and_5958_nl;
  wire[6:0] and_nl;
  wire or_7335_nl;
  wire[1:0] Product2_1_jj_Product2_1_jj_and_1_nl;
  wire[1:0] Product2_1_jj_mux_1_nl;
  wire not_568_nl;
  wire[6:0] Product2_jj_Product2_jj_and_1_nl;
  wire[7:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[16:0] operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[1:0] Product1_mux_3_nl;
  wire[3:0] nnet_linear_layer5_t_result_t_linear_config6_for_mux_5_nl;
  wire or_7367_nl;
  wire[6:0] nnet_linear_layer2_t_layer3_t_linear_config3_for_mux1h_1_nl;
  wire or_7368_nl;
  wire[19:0] mul_nl;
  wire signed [20:0] nl_mul_nl;
  wire[4:0] nnet_product_mult_input_t_config2_weight_t_product_mux_2_nl;
  wire[15:0] nnet_product_mult_input_t_config2_weight_t_product_mux_3_nl;
  wire[15:0] Accum2_mux_133_nl;
  wire[15:0] Accum2_mux_134_nl;
  wire[15:0] Accum2_mux_135_nl;
  wire[15:0] Accum2_1_mux_7_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [47:0] nl_layer6_out_rsci_idat;
  assign nl_layer6_out_rsci_idat = {layer6_out_rsci_idat_47_32 , layer6_out_rsci_idat_31_16
      , layer6_out_rsci_idat_15_0};
  wire [10:0] nl_U_ROM_1i11_1o5_815f6a3dbd0daa2d77beb65dd6cecbbc31_rg_I_1;
  assign nl_U_ROM_1i11_1o5_815f6a3dbd0daa2d77beb65dd6cecbbc31_rg_I_1 = {Accum1_ii_3_0_sva
      , (Result_ires_7_0_sva_1[6:0])};
  wire [8:0] nl_U_ROM_1i9_1o5_4a143e9cb1f27bd26e0331874cec74ad2f_rg_I_1;
  assign nl_U_ROM_1i9_1o5_4a143e9cb1f27bd26e0331874cec74ad2f_rg_I_1 = {z_out_4_8_1
      , (Product2_1_index_acc_sdt[0])};
  wire  nl_myproject_core_core_fsm_inst_Product2_C_0_tr0;
  assign nl_myproject_core_core_fsm_inst_Product2_C_0_tr0 = z_out_2[7];
  wire  nl_myproject_core_core_fsm_inst_Product1_C_1_tr0;
  assign nl_myproject_core_core_fsm_inst_Product1_C_1_tr0 = ~ (z_out_1[3]);
  wire  nl_myproject_core_core_fsm_inst_Accum2_C_0_tr0;
  assign nl_myproject_core_core_fsm_inst_Accum2_C_0_tr0 = z_out_2[7];
  wire  nl_myproject_core_core_fsm_inst_Accum1_C_0_tr0;
  assign nl_myproject_core_core_fsm_inst_Accum1_C_0_tr0 = ~ (z_out_1[3]);
  wire  nl_myproject_core_core_fsm_inst_Product2_1_C_0_tr0;
  assign nl_myproject_core_core_fsm_inst_Product2_1_C_0_tr0 = ~ (z_out_2[2]);
  wire  nl_myproject_core_core_fsm_inst_Accum2_1_C_0_tr0;
  assign nl_myproject_core_core_fsm_inst_Accum2_1_C_0_tr0 = ~ (z_out_2[2]);
  wire  nl_myproject_core_core_fsm_inst_Accum1_1_C_0_tr0;
  assign nl_myproject_core_core_fsm_inst_Accum1_1_C_0_tr0 = z_out_2[7];
  converterBlock_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd224)) input_1_rsci (
      .dat(input_1_rsc_dat),
      .idat(input_1_rsci_idat)
    );
  converterBlock_ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd48)) layer6_out_rsci (
      .idat(nl_layer6_out_rsci_idat[47:0]),
      .dat(layer6_out_rsc_dat)
    );
  converterBlock_ROM_1i11_1o5_4ed11b0fc67dff9823222c14315e503abd  U_ROM_1i11_1o5_815f6a3dbd0daa2d77beb65dd6cecbbc31_rg
      (
      .I_1(nl_U_ROM_1i11_1o5_815f6a3dbd0daa2d77beb65dd6cecbbc31_rg_I_1[10:0]),
      .O_1(ROM_1i11_1o5_815f6a3dbd0daa2d77beb65dd6cecbbc31_1)
    );
  converterBlock_ROM_1i9_1o5_e071483337062336669c4105b16859e3bb  U_ROM_1i9_1o5_4a143e9cb1f27bd26e0331874cec74ad2f_rg
      (
      .I_1(nl_U_ROM_1i9_1o5_4a143e9cb1f27bd26e0331874cec74ad2f_rg_I_1[8:0]),
      .O_1(ROM_1i9_1o5_4a143e9cb1f27bd26e0331874cec74ad2f_1)
    );
  converterBlock_myproject_core_core_fsm myproject_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .Product2_C_0_tr0(nl_myproject_core_core_fsm_inst_Product2_C_0_tr0),
      .Product1_C_1_tr0(nl_myproject_core_core_fsm_inst_Product1_C_1_tr0),
      .Accum2_C_0_tr0(nl_myproject_core_core_fsm_inst_Accum2_C_0_tr0),
      .Accum1_C_0_tr0(nl_myproject_core_core_fsm_inst_Accum1_C_0_tr0),
      .Product2_1_C_0_tr0(nl_myproject_core_core_fsm_inst_Product2_1_C_0_tr0),
      .Result_C_3_tr0(Result_and_1_tmp),
      .Accum2_1_C_0_tr0(nl_myproject_core_core_fsm_inst_Accum2_1_C_0_tr0),
      .Accum1_1_C_0_tr0(nl_myproject_core_core_fsm_inst_Accum1_1_C_0_tr0),
      .Result_1_C_1_tr0(Result_1_Result_1_nor_itm)
    );
  assign and_5052_rgt = and_dcpl_24 & and_dcpl_21 & (fsm_output[4]);
  assign or_6921_rgt = and_5035_cse | (fsm_output[0]);
  assign and_5057_rgt = (Accum1_ii_3_0_sva[1:0]==2'b00) & (fsm_output[11]);
  assign and_5081_rgt = and_dcpl_24 & and_dcpl_41 & (fsm_output[4]);
  assign and_5086_rgt = (Accum1_ii_3_0_sva[1:0]==2'b01) & (fsm_output[11]);
  assign and_5214_rgt = and_dcpl_52 & and_dcpl_60 & (fsm_output[4]);
  assign and_5219_rgt = (Accum1_ii_3_0_sva[1:0]==2'b10) & (fsm_output[11]);
  assign not_2388_nl = ~ (fsm_output[3]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse
      = MUX_v_16_2_2(16'b0000000000000000, z_out_6, not_2388_nl);
  assign Product1_1_ii_or_cse = (fsm_output[5]) | (fsm_output[10]);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_or_cse = Product1_1_ii_or_cse
      | (fsm_output[6]);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 = (Accum2_mux_131[14:10]!=5'b00000);
  assign Accum2_mux_131 = MUX_v_16_128_2(nnet_dense_latency_input_t_layer2_t_config2_acc_0_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_1_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_2_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_3_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_4_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_5_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_6_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_7_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_8_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_9_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_10_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_11_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_12_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_13_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_14_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_15_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_16_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_17_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_18_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_19_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_20_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_21_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_22_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_23_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_24_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_25_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_26_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_27_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_28_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_29_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_30_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_31_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_32_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_33_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_34_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_35_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_36_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_37_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_38_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_39_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_40_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_41_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_42_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_43_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_44_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_45_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_46_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_47_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_48_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_49_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_50_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_51_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_52_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_53_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_54_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_55_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_56_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_57_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_58_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_59_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_60_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_61_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_62_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_63_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_64_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_65_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_66_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_67_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_68_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_69_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_70_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_71_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_72_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_73_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_74_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_75_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_76_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_77_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_78_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_79_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_80_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_81_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_82_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_83_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_84_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_85_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_86_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_87_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_88_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_89_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_90_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_91_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_92_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_93_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_94_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_95_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_96_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_97_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_98_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_99_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_100_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_101_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_102_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_103_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_104_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_105_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_106_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_107_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_108_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_109_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_110_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_111_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_112_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_113_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_114_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_115_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_116_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_117_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_118_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_119_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_120_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_121_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_122_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_123_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_124_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_125_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_126_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_127_lpi_3, Result_ires_7_0_sva_1[6:0]);
  assign operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl =  -conv_s2s_16_17(Accum2_mux_131);
  assign operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1 = readslicef_17_1_16(operator_16_6_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign Accum2_1_mux_6 = MUX_v_16_3_2(nnet_dense_latency_input_t_layer2_t_config2_acc_0_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_acc_1_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_acc_10_lpi_3,
      Accum1_ii_3_0_sva[1:0]);
  assign Result_and_1_tmp = (Result_ires_7_0_sva_1[7]) & (nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[7])
      & (nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_7_0_sva_1[7]) & (z_out_2[7]);
  assign or_dcpl_69 = (Accum1_ii_3_0_sva[1:0]!=2'b01);
  assign or_dcpl_70 = or_dcpl_69 | (~ (Accum1_ii_3_0_sva[3]));
  assign or_dcpl_80 = (Accum1_ii_3_0_sva[1:0]!=2'b00);
  assign or_dcpl_81 = or_dcpl_80 | (Accum1_ii_3_0_sva[3]);
  assign or_dcpl_420 = or_dcpl_80 | (~ (Accum1_ii_3_0_sva[3]));
  assign or_dcpl_423 = or_dcpl_69 | (Accum1_ii_3_0_sva[3]);
  assign or_dcpl_682 = ~((Accum1_ii_3_0_sva[1:0]==2'b11));
  assign or_dcpl_683 = or_dcpl_682 | (~ (Accum1_ii_3_0_sva[3]));
  assign or_dcpl_686 = (Accum1_ii_3_0_sva[1:0]!=2'b10);
  assign or_dcpl_687 = or_dcpl_686 | (Accum1_ii_3_0_sva[3]);
  assign or_dcpl_946 = or_dcpl_686 | (~ (Accum1_ii_3_0_sva[3]));
  assign or_dcpl_949 = or_dcpl_682 | (Accum1_ii_3_0_sva[3]);
  assign and_dcpl_2 = ~((fsm_output[14:13]!=2'b00));
  assign or_dcpl_2015 = (nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[1:0]!=2'b01);
  assign or_dcpl_2016 = (nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[1:0]!=2'b10);
  assign or_dcpl_2020 = (fsm_output[14:13]!=2'b00);
  assign or_dcpl_2027 = (Result_ires_7_0_sva_1[3:2]!=2'b00);
  assign or_dcpl_2028 = (Result_ires_7_0_sva_1[6]) | (Result_ires_7_0_sva_1[1]);
  assign or_dcpl_2029 = or_dcpl_2028 | (Result_ires_7_0_sva_1[0]);
  assign or_dcpl_2030 = or_dcpl_2029 | or_dcpl_2027;
  assign or_dcpl_2031 = (Accum1_ii_3_0_sva[2]) | (Result_ires_7_0_sva_1[4]);
  assign or_dcpl_2032 = or_dcpl_2031 | (Result_ires_7_0_sva_1[5]);
  assign or_dcpl_2035 = or_dcpl_81 | or_dcpl_2032;
  assign or_dcpl_2037 = or_dcpl_2028 | (~ (Result_ires_7_0_sva_1[0]));
  assign or_dcpl_2038 = or_dcpl_2037 | or_dcpl_2027;
  assign or_dcpl_2040 = (Result_ires_7_0_sva_1[3:2]!=2'b10);
  assign or_dcpl_2041 = (Result_ires_7_0_sva_1[6]) | (~ (Result_ires_7_0_sva_1[1]));
  assign or_dcpl_2042 = or_dcpl_2041 | (Result_ires_7_0_sva_1[0]);
  assign or_dcpl_2043 = or_dcpl_2042 | or_dcpl_2040;
  assign or_dcpl_2045 = (Result_ires_7_0_sva_1[3:2]!=2'b01);
  assign or_dcpl_2046 = (~ (Result_ires_7_0_sva_1[6])) | (Result_ires_7_0_sva_1[1]);
  assign or_dcpl_2047 = or_dcpl_2046 | (Result_ires_7_0_sva_1[0]);
  assign or_dcpl_2048 = or_dcpl_2047 | or_dcpl_2045;
  assign or_dcpl_2049 = or_dcpl_2031 | (~ (Result_ires_7_0_sva_1[5]));
  assign or_dcpl_2050 = or_dcpl_81 | or_dcpl_2049;
  assign or_dcpl_2052 = or_dcpl_2047 | or_dcpl_2040;
  assign or_dcpl_2053 = (~ (Accum1_ii_3_0_sva[2])) | (Result_ires_7_0_sva_1[4]);
  assign or_dcpl_2054 = or_dcpl_2053 | (~ (Result_ires_7_0_sva_1[5]));
  assign or_dcpl_2057 = or_dcpl_949 | or_dcpl_2054;
  assign or_dcpl_2059 = or_dcpl_2046 | (~ (Result_ires_7_0_sva_1[0]));
  assign or_dcpl_2060 = or_dcpl_2059 | or_dcpl_2040;
  assign or_dcpl_2062 = ~((Result_ires_7_0_sva_1[6]) & (Result_ires_7_0_sva_1[1]));
  assign or_dcpl_2063 = or_dcpl_2062 | (Result_ires_7_0_sva_1[0]);
  assign or_dcpl_2064 = or_dcpl_2063 | or_dcpl_2040;
  assign or_dcpl_2066 = or_dcpl_2062 | (~ (Result_ires_7_0_sva_1[0]));
  assign or_dcpl_2067 = or_dcpl_2066 | or_dcpl_2040;
  assign or_dcpl_2069 = ~((Result_ires_7_0_sva_1[3:2]==2'b11));
  assign or_dcpl_2070 = or_dcpl_2047 | or_dcpl_2069;
  assign or_dcpl_2072 = or_dcpl_2059 | or_dcpl_2069;
  assign or_dcpl_2074 = or_dcpl_2063 | or_dcpl_2069;
  assign or_dcpl_2076 = or_dcpl_2066 | or_dcpl_2069;
  assign or_dcpl_2078 = or_dcpl_2047 | or_dcpl_2027;
  assign or_dcpl_2079 = ~((Accum1_ii_3_0_sva[2]) & (Result_ires_7_0_sva_1[4]));
  assign or_dcpl_2080 = or_dcpl_2079 | (~ (Result_ires_7_0_sva_1[5]));
  assign or_dcpl_2081 = or_dcpl_949 | or_dcpl_2080;
  assign or_dcpl_2083 = or_dcpl_2059 | or_dcpl_2027;
  assign or_dcpl_2085 = or_dcpl_2059 | or_dcpl_2045;
  assign or_dcpl_2087 = or_dcpl_2063 | or_dcpl_2027;
  assign or_dcpl_2089 = or_dcpl_2066 | or_dcpl_2027;
  assign or_dcpl_2093 = or_dcpl_2063 | or_dcpl_2045;
  assign or_dcpl_2095 = or_dcpl_2066 | or_dcpl_2045;
  assign or_dcpl_2107 = or_dcpl_420 | or_dcpl_2032;
  assign or_dcpl_2110 = or_dcpl_2042 | or_dcpl_2027;
  assign or_dcpl_2112 = or_dcpl_2041 | (~ (Result_ires_7_0_sva_1[0]));
  assign or_dcpl_2113 = or_dcpl_2112 | or_dcpl_2027;
  assign or_dcpl_2115 = or_dcpl_2029 | or_dcpl_2045;
  assign or_dcpl_2117 = or_dcpl_2037 | or_dcpl_2045;
  assign or_dcpl_2120 = or_dcpl_2042 | or_dcpl_2045;
  assign or_dcpl_2122 = or_dcpl_2112 | or_dcpl_2045;
  assign or_dcpl_2124 = or_dcpl_2029 | or_dcpl_2040;
  assign or_dcpl_2126 = or_dcpl_2037 | or_dcpl_2040;
  assign or_dcpl_2129 = or_dcpl_2112 | or_dcpl_2040;
  assign or_dcpl_2131 = or_dcpl_2029 | or_dcpl_2069;
  assign or_dcpl_2133 = or_dcpl_2037 | or_dcpl_2069;
  assign or_dcpl_2135 = or_dcpl_2042 | or_dcpl_2069;
  assign or_dcpl_2137 = or_dcpl_2112 | or_dcpl_2069;
  assign or_dcpl_2140 = (Accum1_ii_3_0_sva[2]) | (~ (Result_ires_7_0_sva_1[4]));
  assign or_dcpl_2141 = or_dcpl_2140 | (Result_ires_7_0_sva_1[5]);
  assign or_dcpl_2142 = or_dcpl_420 | or_dcpl_2141;
  assign or_dcpl_2160 = or_dcpl_420 | or_dcpl_2049;
  assign or_dcpl_2179 = or_dcpl_2140 | (~ (Result_ires_7_0_sva_1[5]));
  assign or_dcpl_2180 = or_dcpl_420 | or_dcpl_2179;
  assign or_dcpl_2234 = or_dcpl_81 | or_dcpl_2179;
  assign or_dcpl_2273 = or_dcpl_70 | or_dcpl_2032;
  assign or_dcpl_2291 = or_dcpl_70 | or_dcpl_2141;
  assign or_dcpl_2310 = or_dcpl_70 | or_dcpl_2049;
  assign or_dcpl_2330 = or_dcpl_70 | or_dcpl_2179;
  assign or_dcpl_2419 = or_dcpl_423 | or_dcpl_2032;
  assign or_dcpl_2423 = or_dcpl_946 | or_dcpl_2032;
  assign or_dcpl_2441 = or_dcpl_946 | or_dcpl_2141;
  assign or_dcpl_2461 = or_dcpl_946 | or_dcpl_2049;
  assign or_dcpl_2479 = or_dcpl_946 | or_dcpl_2179;
  assign or_dcpl_2570 = or_dcpl_683 | or_dcpl_2032;
  assign or_dcpl_2589 = or_dcpl_683 | or_dcpl_2141;
  assign or_dcpl_2607 = or_dcpl_423 | or_dcpl_2141;
  assign or_dcpl_2609 = or_dcpl_683 | or_dcpl_2049;
  assign or_dcpl_2627 = or_dcpl_683 | or_dcpl_2179;
  assign or_dcpl_2717 = or_dcpl_2053 | (Result_ires_7_0_sva_1[5]);
  assign or_dcpl_2718 = or_dcpl_420 | or_dcpl_2717;
  assign or_dcpl_2737 = or_dcpl_2079 | (Result_ires_7_0_sva_1[5]);
  assign or_dcpl_2738 = or_dcpl_420 | or_dcpl_2737;
  assign or_dcpl_2756 = or_dcpl_420 | or_dcpl_2054;
  assign or_dcpl_2775 = or_dcpl_420 | or_dcpl_2080;
  assign or_dcpl_2793 = or_dcpl_81 | or_dcpl_2141;
  assign or_dcpl_2795 = or_dcpl_423 | or_dcpl_2049;
  assign or_dcpl_2867 = or_dcpl_70 | or_dcpl_2717;
  assign or_dcpl_2886 = or_dcpl_70 | or_dcpl_2737;
  assign or_dcpl_2904 = or_dcpl_70 | or_dcpl_2054;
  assign or_dcpl_2924 = or_dcpl_70 | or_dcpl_2080;
  assign or_dcpl_2977 = or_dcpl_423 | or_dcpl_2179;
  assign or_dcpl_3100 = or_dcpl_687 | or_dcpl_2032;
  assign or_dcpl_3119 = or_dcpl_687 | or_dcpl_2141;
  assign or_dcpl_3137 = or_dcpl_687 | or_dcpl_2049;
  assign or_dcpl_3157 = or_dcpl_687 | or_dcpl_2179;
  assign or_dcpl_3246 = or_dcpl_949 | or_dcpl_2032;
  assign or_dcpl_3266 = or_dcpl_949 | or_dcpl_2141;
  assign or_dcpl_3284 = or_dcpl_949 | or_dcpl_2049;
  assign or_dcpl_3303 = or_dcpl_949 | or_dcpl_2179;
  assign or_dcpl_3393 = or_dcpl_81 | or_dcpl_2717;
  assign or_dcpl_3411 = or_dcpl_81 | or_dcpl_2737;
  assign or_dcpl_3430 = or_dcpl_81 | or_dcpl_2054;
  assign or_dcpl_3449 = or_dcpl_81 | or_dcpl_2080;
  assign or_dcpl_3539 = or_dcpl_423 | or_dcpl_2717;
  assign or_dcpl_3557 = or_dcpl_423 | or_dcpl_2737;
  assign or_dcpl_3576 = or_dcpl_423 | or_dcpl_2054;
  assign or_dcpl_3594 = or_dcpl_423 | or_dcpl_2080;
  assign or_dcpl_3684 = or_dcpl_687 | or_dcpl_2717;
  assign or_dcpl_3703 = or_dcpl_687 | or_dcpl_2737;
  assign or_dcpl_3723 = or_dcpl_687 | or_dcpl_2054;
  assign or_dcpl_3741 = or_dcpl_687 | or_dcpl_2080;
  assign or_dcpl_3830 = or_dcpl_949 | or_dcpl_2717;
  assign or_dcpl_3850 = or_dcpl_949 | or_dcpl_2737;
  assign or_dcpl_3947 = (z_out_4_8_1[5]) | (Product2_1_index_acc_sdt[0]);
  assign or_dcpl_3948 = (z_out_4_8_1[4:3]!=2'b00);
  assign or_dcpl_3949 = or_dcpl_3948 | or_dcpl_3947;
  assign or_dcpl_3950 = (z_out_4_8_1[2:1]!=2'b00);
  assign or_dcpl_3951 = (z_out_4_8_1[7:6]!=2'b00);
  assign or_dcpl_3952 = or_dcpl_3951 | (z_out_4_8_1[0]);
  assign or_dcpl_3953 = or_dcpl_3952 | or_dcpl_3950;
  assign or_dcpl_3955 = (z_out_4_8_1[5]) | (~ (Product2_1_index_acc_sdt[0]));
  assign or_dcpl_3956 = or_dcpl_3948 | or_dcpl_3955;
  assign or_dcpl_3958 = (z_out_4_8_1[2:1]!=2'b10);
  assign or_dcpl_3959 = or_dcpl_3951 | (~ (z_out_4_8_1[0]));
  assign or_dcpl_3960 = or_dcpl_3959 | or_dcpl_3958;
  assign or_dcpl_3962 = (~ (z_out_4_8_1[5])) | (Product2_1_index_acc_sdt[0]);
  assign or_dcpl_3963 = (z_out_4_8_1[4:3]!=2'b10);
  assign or_dcpl_3964 = or_dcpl_3963 | or_dcpl_3962;
  assign or_dcpl_3965 = (z_out_4_8_1[2:1]!=2'b01);
  assign or_dcpl_3966 = or_dcpl_3952 | or_dcpl_3965;
  assign or_dcpl_3968 = ~((z_out_4_8_1[5]) & (Product2_1_index_acc_sdt[0]));
  assign or_dcpl_3969 = or_dcpl_3963 | or_dcpl_3968;
  assign or_dcpl_3971 = or_dcpl_3959 | or_dcpl_3965;
  assign or_dcpl_3974 = or_dcpl_3952 | or_dcpl_3958;
  assign or_dcpl_3979 = ~((z_out_4_8_1[2:1]==2'b11));
  assign or_dcpl_3980 = or_dcpl_3952 | or_dcpl_3979;
  assign or_dcpl_3984 = or_dcpl_3959 | or_dcpl_3979;
  assign or_dcpl_3987 = ~((z_out_4_8_1[4:3]==2'b11));
  assign or_dcpl_3988 = or_dcpl_3987 | or_dcpl_3962;
  assign or_dcpl_3990 = or_dcpl_3987 | or_dcpl_3968;
  assign or_dcpl_3992 = or_dcpl_3959 | or_dcpl_3950;
  assign or_dcpl_4008 = (z_out_4_8_1[7:6]!=2'b01);
  assign or_dcpl_4009 = or_dcpl_4008 | (z_out_4_8_1[0]);
  assign or_dcpl_4010 = or_dcpl_4009 | or_dcpl_3950;
  assign or_dcpl_4014 = or_dcpl_4008 | (~ (z_out_4_8_1[0]));
  assign or_dcpl_4015 = or_dcpl_4014 | or_dcpl_3950;
  assign or_dcpl_4018 = or_dcpl_4009 | or_dcpl_3965;
  assign or_dcpl_4021 = or_dcpl_4014 | or_dcpl_3965;
  assign or_dcpl_4024 = or_dcpl_4009 | or_dcpl_3958;
  assign or_dcpl_4027 = or_dcpl_4014 | or_dcpl_3958;
  assign or_dcpl_4031 = or_dcpl_4009 | or_dcpl_3979;
  assign or_dcpl_4034 = or_dcpl_4014 | or_dcpl_3979;
  assign or_dcpl_4037 = (z_out_4_8_1[4:3]!=2'b01);
  assign or_dcpl_4038 = or_dcpl_4037 | or_dcpl_3947;
  assign or_dcpl_4040 = or_dcpl_4037 | or_dcpl_3955;
  assign or_dcpl_4058 = or_dcpl_3963 | or_dcpl_3947;
  assign or_dcpl_4060 = or_dcpl_3963 | or_dcpl_3955;
  assign or_dcpl_4077 = or_dcpl_3987 | or_dcpl_3947;
  assign or_dcpl_4079 = or_dcpl_3987 | or_dcpl_3955;
  assign or_dcpl_4097 = or_dcpl_3948 | or_dcpl_3962;
  assign or_dcpl_4099 = or_dcpl_3948 | or_dcpl_3968;
  assign or_dcpl_4117 = or_dcpl_4037 | or_dcpl_3962;
  assign or_dcpl_4119 = or_dcpl_4037 | or_dcpl_3968;
  assign or_dcpl_4172 = (z_out_4_8_1[7:6]!=2'b10);
  assign or_dcpl_4173 = or_dcpl_4172 | (z_out_4_8_1[0]);
  assign or_dcpl_4174 = or_dcpl_4173 | or_dcpl_3950;
  assign or_dcpl_4177 = or_dcpl_4172 | (~ (z_out_4_8_1[0]));
  assign or_dcpl_4178 = or_dcpl_4177 | or_dcpl_3950;
  assign or_dcpl_4182 = or_dcpl_4173 | or_dcpl_3965;
  assign or_dcpl_4185 = or_dcpl_4177 | or_dcpl_3965;
  assign or_dcpl_4188 = or_dcpl_4173 | or_dcpl_3958;
  assign or_dcpl_4191 = or_dcpl_4177 | or_dcpl_3958;
  assign or_dcpl_4194 = or_dcpl_4173 | or_dcpl_3979;
  assign or_dcpl_4198 = or_dcpl_4177 | or_dcpl_3979;
  assign or_dcpl_4396 = (Result_ires_7_0_sva_1[0]) | (Result_ires_7_0_sva_1[2]);
  assign or_dcpl_4397 = or_dcpl_4396 | (Result_ires_7_0_sva_1[3]);
  assign or_dcpl_4398 = (Result_ires_7_0_sva_1[5:4]!=2'b00);
  assign or_dcpl_4399 = or_dcpl_4398 | or_dcpl_2028;
  assign and_dcpl_20 = ~((Result_ires_7_0_sva_1[0]) | (Result_ires_7_0_sva_1[2]));
  assign and_dcpl_21 = and_dcpl_20 & (~ (Result_ires_7_0_sva_1[3]));
  assign and_dcpl_22 = ~((Result_ires_7_0_sva_1[6]) | (Result_ires_7_0_sva_1[1]));
  assign and_dcpl_23 = ~((Result_ires_7_0_sva_1[5:4]!=2'b00));
  assign and_dcpl_24 = and_dcpl_23 & and_dcpl_22;
  assign and_dcpl_31 = (Result_ires_7_0_sva_1[0]) & (Result_ires_7_0_sva_1[2]);
  assign and_dcpl_32 = and_dcpl_31 & (Result_ires_7_0_sva_1[3]);
  assign and_dcpl_33 = (Result_ires_7_0_sva_1[6]) & (Result_ires_7_0_sva_1[1]);
  assign and_dcpl_34 = (Result_ires_7_0_sva_1[5:4]==2'b11);
  assign and_dcpl_35 = and_dcpl_34 & and_dcpl_33;
  assign or_dcpl_4409 = ~((Result_ires_7_0_sva_1[0]) & (Result_ires_7_0_sva_1[2]));
  assign or_dcpl_4410 = or_dcpl_4409 | (~ (Result_ires_7_0_sva_1[3]));
  assign or_dcpl_4411 = ~((Result_ires_7_0_sva_1[5:4]==2'b11));
  assign or_dcpl_4412 = or_dcpl_4411 | or_dcpl_2062;
  assign and_dcpl_37 = (~ (Result_ires_7_0_sva_1[0])) & (Result_ires_7_0_sva_1[2]);
  assign and_dcpl_38 = and_dcpl_37 & (Result_ires_7_0_sva_1[3]);
  assign or_dcpl_4414 = (Result_ires_7_0_sva_1[0]) | (~ (Result_ires_7_0_sva_1[2]));
  assign or_dcpl_4415 = or_dcpl_4414 | (~ (Result_ires_7_0_sva_1[3]));
  assign and_dcpl_40 = (Result_ires_7_0_sva_1[0]) & (~ (Result_ires_7_0_sva_1[2]));
  assign and_dcpl_41 = and_dcpl_40 & (~ (Result_ires_7_0_sva_1[3]));
  assign or_dcpl_4419 = (~ (Result_ires_7_0_sva_1[0])) | (Result_ires_7_0_sva_1[2]);
  assign or_dcpl_4420 = or_dcpl_4419 | (Result_ires_7_0_sva_1[3]);
  assign and_dcpl_48 = (Result_ires_7_0_sva_1[6]) & (~ (Result_ires_7_0_sva_1[1]));
  assign and_dcpl_49 = and_dcpl_34 & and_dcpl_48;
  assign or_dcpl_4422 = or_dcpl_4411 | or_dcpl_2046;
  assign and_dcpl_51 = (~ (Result_ires_7_0_sva_1[6])) & (Result_ires_7_0_sva_1[1]);
  assign and_dcpl_52 = and_dcpl_23 & and_dcpl_51;
  assign or_dcpl_4424 = or_dcpl_4398 | or_dcpl_2041;
  assign and_dcpl_56 = and_dcpl_40 & (Result_ires_7_0_sva_1[3]);
  assign or_dcpl_4428 = or_dcpl_4419 | (~ (Result_ires_7_0_sva_1[3]));
  assign and_dcpl_58 = and_dcpl_37 & (~ (Result_ires_7_0_sva_1[3]));
  assign or_dcpl_4430 = or_dcpl_4414 | (Result_ires_7_0_sva_1[3]);
  assign and_dcpl_60 = and_dcpl_20 & (Result_ires_7_0_sva_1[3]);
  assign or_dcpl_4432 = or_dcpl_4396 | (~ (Result_ires_7_0_sva_1[3]));
  assign and_dcpl_62 = and_dcpl_31 & (~ (Result_ires_7_0_sva_1[3]));
  assign or_dcpl_4434 = or_dcpl_4409 | (Result_ires_7_0_sva_1[3]);
  assign and_dcpl_85 = (Result_ires_7_0_sva_1[5:4]==2'b10);
  assign and_dcpl_86 = and_dcpl_85 & and_dcpl_33;
  assign or_dcpl_4456 = (Result_ires_7_0_sva_1[5:4]!=2'b10);
  assign or_dcpl_4457 = or_dcpl_4456 | or_dcpl_2062;
  assign and_dcpl_88 = (Result_ires_7_0_sva_1[5:4]==2'b01);
  assign and_dcpl_89 = and_dcpl_88 & and_dcpl_22;
  assign or_dcpl_4459 = (Result_ires_7_0_sva_1[5:4]!=2'b01);
  assign or_dcpl_4460 = or_dcpl_4459 | or_dcpl_2028;
  assign and_dcpl_93 = and_dcpl_85 & and_dcpl_48;
  assign or_dcpl_4464 = or_dcpl_4456 | or_dcpl_2046;
  assign and_dcpl_95 = and_dcpl_88 & and_dcpl_51;
  assign or_dcpl_4466 = or_dcpl_4459 | or_dcpl_2041;
  assign and_dcpl_123 = and_dcpl_88 & and_dcpl_33;
  assign or_dcpl_4494 = or_dcpl_4459 | or_dcpl_2062;
  assign and_dcpl_125 = and_dcpl_85 & and_dcpl_22;
  assign or_dcpl_4496 = or_dcpl_4456 | or_dcpl_2028;
  assign and_dcpl_129 = and_dcpl_88 & and_dcpl_48;
  assign or_dcpl_4500 = or_dcpl_4459 | or_dcpl_2046;
  assign and_dcpl_131 = and_dcpl_85 & and_dcpl_51;
  assign or_dcpl_4502 = or_dcpl_4456 | or_dcpl_2041;
  assign and_dcpl_159 = and_dcpl_23 & and_dcpl_33;
  assign or_dcpl_4530 = or_dcpl_4398 | or_dcpl_2062;
  assign and_dcpl_161 = and_dcpl_34 & and_dcpl_22;
  assign or_dcpl_4532 = or_dcpl_4411 | or_dcpl_2028;
  assign and_dcpl_165 = and_dcpl_23 & and_dcpl_48;
  assign or_dcpl_4536 = or_dcpl_4398 | or_dcpl_2046;
  assign and_dcpl_167 = and_dcpl_34 & and_dcpl_51;
  assign or_dcpl_4538 = or_dcpl_4411 | or_dcpl_2041;
  assign and_5035_cse = Result_and_1_tmp & (fsm_output[10]);
  assign and_5068_cse = (fsm_output[10:5]!=6'b000000);
  assign or_tmp_2362 = (fsm_output[2:0]!=3'b000) | and_5035_cse;
  assign or_tmp_2754 = (fsm_output[9:7]!=3'b000);
  assign Accum1_ii_3_0_sva_mx0c0 = ((~ (z_out_1[3])) & (fsm_output[3])) | (fsm_output[0]);
  assign Accum1_ii_3_0_sva_mx0c3 = or_dcpl_2020 | (fsm_output[12:8]!=5'b00000);
  assign nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1_mx0c2 = or_dcpl_2020
      | (fsm_output[12]);
  assign Product2_1_index_mux_cse = MUX_v_7_2_2(Product1_1_ii_7_0_sva_6_0, (Result_ires_7_0_sva_1[6:0]),
      fsm_output[11]);
  assign or_7342_cse = (fsm_output[13]) | (fsm_output[11]) | (fsm_output[9]);
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_31_16_lpi_2
          <= 16'b0000000000000000;
    end
    else if ( (~ or_dcpl_2015) & (fsm_output[13]) ) begin
      nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_31_16_lpi_2
          <= Accum2_1_mux_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_47_32_lpi_2
          <= 16'b0000000000000000;
    end
    else if ( (~ or_dcpl_2016) & (fsm_output[13]) ) begin
      nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_47_32_lpi_2
          <= Accum2_1_mux_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer6_out_rsci_idat_15_0 <= 16'b0000000000000000;
    end
    else if ( fsm_output[13] ) begin
      layer6_out_rsci_idat_15_0 <= MUX_v_16_2_2(nnet_dense_latency_input_t_layer2_t_config2_acc_100_lpi_3,
          Accum2_1_mux_6, and_655_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer6_out_rsci_idat_31_16 <= 16'b0000000000000000;
    end
    else if ( fsm_output[13] ) begin
      layer6_out_rsci_idat_31_16 <= MUX_v_16_2_2(Accum2_1_mux_6, nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_31_16_lpi_2,
          and_661_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer6_out_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else if ( fsm_output[13] ) begin
      layer6_out_rsci_idat_47_32 <= MUX_v_16_2_2(Accum2_1_mux_6, nnet_linear_layer5_t_result_t_linear_config6_for_io_read_layer6_out_rsc_sdt_47_32_lpi_2,
          and_667_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Accum1_ii_3_0_sva <= 4'b0000;
    end
    else if ( Accum1_ii_3_0_sva_mx0c0 | ((z_out_1[3]) & (fsm_output[3])) | (fsm_output[5])
        | Accum1_ii_3_0_sva_mx0c3 ) begin
      Accum1_ii_3_0_sva <= MUX_v_4_2_2(4'b0000, Product1_ii_Product1_ii_mux_nl, Accum1_ii_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_0_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_0_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_10_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_10_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_100_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_100_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1000_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1000_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1001_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1001_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1002_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1002_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1003_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1003_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1004_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1004_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1005_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1005_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1006_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1006_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1007_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1007_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1008_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1008_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1009_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1009_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_101_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_101_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1010_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1010_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1011_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1011_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1012_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1012_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1013_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1013_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1014_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1014_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1015_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1015_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1016_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1016_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1017_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1017_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1018_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1018_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1019_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1019_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_102_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_102_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1020_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1020_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1021_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1021_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1022_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1022_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1023_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1023_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1024_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_2107 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1024_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1025_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1025_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1026_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1026_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1027_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1027_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1028_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1028_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1029_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1029_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_103_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_103_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1030_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1030_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1031_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1031_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1032_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1032_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1033_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1033_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1034_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1034_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1035_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1035_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1036_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1036_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1037_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1037_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1038_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1038_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1039_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1039_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_104_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_104_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1040_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1040_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1041_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1041_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1042_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1042_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1043_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1043_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1044_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1044_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1045_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1045_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1046_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1046_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1047_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1047_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1048_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1048_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1049_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1049_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_105_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_105_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1050_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1050_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1051_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1051_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1052_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1052_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1053_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1053_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1054_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1054_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1055_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1055_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1056_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1056_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1057_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1057_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1058_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1058_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1059_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1059_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_106_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_106_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1060_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1060_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1061_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1061_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1062_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1062_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1063_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1063_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1064_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1064_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1065_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1065_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1066_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1066_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1067_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1067_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1068_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1068_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1069_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1069_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_107_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_107_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1070_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1070_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1071_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1071_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1072_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1072_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1073_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1073_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1074_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1074_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1075_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1075_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1076_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1076_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1077_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1077_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1078_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1078_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1079_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1079_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_108_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_108_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1080_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1080_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1081_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1081_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1082_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1082_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1083_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1083_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1084_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1084_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1085_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1085_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1086_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1086_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1087_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1087_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1088_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1088_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1089_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1089_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_109_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_109_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1090_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1090_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1091_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1091_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1092_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1092_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1093_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1093_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1094_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1094_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1095_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1095_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1096_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1096_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1097_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1097_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1098_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1098_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1099_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1099_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_11_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_11_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_110_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_110_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1100_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1100_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1101_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1101_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1102_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1102_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1103_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2107 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1103_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1104_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1104_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1105_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1105_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1106_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1106_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1107_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1107_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1108_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1108_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1109_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1109_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_111_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_111_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1110_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1110_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1111_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1111_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1112_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1112_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1113_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1113_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1114_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1114_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1115_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1115_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1116_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1116_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1117_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1117_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1118_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1118_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1119_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2142 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1119_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_112_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_112_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1120_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1120_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1121_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1121_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1122_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1122_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1123_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1123_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1124_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1124_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1125_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1125_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1126_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1126_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1127_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1127_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1128_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1128_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1129_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1129_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_113_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_113_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1130_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1130_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1131_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1131_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1132_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1132_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1133_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1133_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1134_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1134_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1135_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2160 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1135_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1136_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1136_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1137_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1137_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1138_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1138_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1139_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1139_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_114_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_114_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1140_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1140_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1141_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1141_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1142_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1142_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1143_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1143_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1144_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1144_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1145_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1145_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1146_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1146_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1147_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1147_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1148_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1148_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1149_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1149_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_115_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_115_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1150_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1150_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1151_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2180 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1151_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1152_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_2273 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1152_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1153_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1153_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1154_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1154_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1155_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1155_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1156_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1156_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1157_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1157_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1158_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1158_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1159_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1159_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_116_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_116_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1160_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1160_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1161_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1161_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1162_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1162_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1163_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1163_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1164_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1164_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1165_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1165_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1166_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1166_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1167_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1167_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1168_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1168_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1169_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1169_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_117_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_117_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1170_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1170_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1171_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1171_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1172_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1172_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1173_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1173_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1174_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1174_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1175_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1175_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1176_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1176_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1177_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1177_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1178_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1178_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1179_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1179_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_118_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_118_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1180_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1180_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1181_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1181_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1182_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1182_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1183_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1183_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1184_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1184_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1185_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1185_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1186_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1186_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1187_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1187_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1188_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1188_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1189_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1189_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_119_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_119_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1190_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1190_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1191_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1191_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1192_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1192_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1193_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1193_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1194_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1194_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1195_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1195_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1196_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1196_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1197_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1197_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1198_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1198_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1199_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1199_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_12_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_12_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_120_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_120_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1200_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1200_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1201_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1201_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1202_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1202_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1203_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1203_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1204_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1204_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1205_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1205_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1206_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1206_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1207_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1207_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1208_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1208_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1209_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1209_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_121_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_121_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1210_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1210_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1211_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1211_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1212_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1212_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1213_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1213_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1214_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1214_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1215_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1215_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1216_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1216_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1217_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1217_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1218_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1218_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1219_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1219_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_122_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_122_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1220_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1220_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1221_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1221_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1222_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1222_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1223_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1223_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1224_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1224_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1225_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1225_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1226_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1226_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1227_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1227_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1228_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1228_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1229_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1229_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_123_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_123_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1230_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1230_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1231_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2273 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1231_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1232_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1232_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1233_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1233_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1234_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1234_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1235_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1235_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1236_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1236_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1237_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1237_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1238_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1238_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1239_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1239_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_124_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_124_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1240_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1240_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1241_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1241_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1242_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1242_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1243_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1243_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1244_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1244_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1245_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1245_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1246_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1246_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1247_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2291 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1247_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1248_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1248_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1249_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1249_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_125_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_125_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1250_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1250_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1251_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1251_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1252_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1252_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1253_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1253_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1254_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1254_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1255_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1255_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1256_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1256_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1257_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1257_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1258_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1258_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1259_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1259_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_126_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_126_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1260_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1260_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1261_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1261_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1262_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1262_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1263_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2310 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1263_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1264_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1264_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1265_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1265_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1266_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1266_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1267_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1267_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1268_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1268_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1269_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1269_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_127_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_127_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1270_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1270_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1271_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1271_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1272_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1272_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1273_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1273_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1274_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1274_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1275_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1275_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1276_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1276_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1277_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1277_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1278_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1278_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1279_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2330 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1279_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_128_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_2419 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_128_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1280_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_2423 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1280_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1281_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1281_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1282_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1282_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1283_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1283_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1284_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1284_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1285_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1285_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1286_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1286_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1287_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1287_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1288_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1288_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1289_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1289_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_129_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_129_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1290_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1290_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1291_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1291_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1292_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1292_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1293_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1293_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1294_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1294_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1295_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1295_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1296_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1296_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1297_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1297_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1298_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1298_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1299_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1299_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_13_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_13_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_130_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_130_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1300_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1300_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1301_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1301_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1302_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1302_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1303_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1303_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1304_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1304_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1305_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1305_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1306_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1306_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1307_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1307_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1308_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1308_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1309_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1309_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_131_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_131_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1310_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1310_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1311_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1311_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1312_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1312_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1313_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1313_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1314_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1314_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1315_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1315_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1316_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1316_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1317_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1317_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1318_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1318_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1319_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1319_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_132_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_132_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1320_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1320_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1321_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1321_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1322_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1322_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1323_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1323_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1324_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1324_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1325_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1325_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1326_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1326_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1327_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1327_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1328_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1328_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1329_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1329_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_133_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_133_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1330_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1330_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1331_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1331_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1332_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1332_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1333_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1333_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1334_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1334_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1335_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1335_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1336_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1336_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1337_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1337_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1338_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1338_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1339_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1339_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_134_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_134_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1340_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1340_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1341_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1341_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1342_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1342_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1343_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1343_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1344_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1344_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1345_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1345_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1346_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1346_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1347_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1347_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1348_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1348_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1349_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1349_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_135_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_135_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1350_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1350_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1351_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1351_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1352_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1352_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1353_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1353_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1354_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1354_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1355_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1355_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1356_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1356_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1357_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1357_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1358_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1358_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1359_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2423 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1359_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_136_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_136_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1360_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1360_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1361_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1361_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1362_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1362_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1363_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1363_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1364_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1364_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1365_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1365_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1366_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1366_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1367_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1367_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1368_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1368_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1369_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1369_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_137_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_137_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1370_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1370_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1371_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1371_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1372_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1372_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1373_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1373_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1374_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1374_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1375_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2441 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1375_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1376_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1376_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1377_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1377_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1378_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1378_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1379_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1379_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_138_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_138_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1380_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1380_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1381_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1381_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1382_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1382_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1383_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1383_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1384_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1384_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1385_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1385_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1386_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1386_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1387_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1387_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1388_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1388_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1389_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1389_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_139_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_139_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1390_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1390_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1391_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2461 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1391_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1392_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1392_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1393_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1393_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1394_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1394_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1395_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1395_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1396_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1396_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1397_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1397_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1398_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1398_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1399_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1399_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_14_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_14_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_140_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_140_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1400_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1400_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1401_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1401_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1402_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1402_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1403_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1403_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1404_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1404_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1405_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1405_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1406_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1406_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1407_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2479 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1407_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1408_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_2570 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1408_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1409_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1409_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_141_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_141_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1410_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1410_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1411_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1411_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1412_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1412_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1413_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1413_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1414_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1414_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1415_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1415_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1416_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1416_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1417_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1417_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1418_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1418_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1419_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1419_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_142_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_142_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1420_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1420_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1421_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1421_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1422_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1422_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1423_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1423_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1424_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1424_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1425_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1425_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1426_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1426_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1427_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1427_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1428_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1428_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1429_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1429_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_143_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_143_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1430_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1430_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1431_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1431_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1432_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1432_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1433_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1433_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1434_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1434_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1435_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1435_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1436_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1436_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1437_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1437_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1438_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1438_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1439_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1439_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_144_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_144_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1440_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1440_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1441_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1441_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1442_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1442_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1443_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1443_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1444_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1444_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1445_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1445_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1446_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1446_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1447_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1447_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1448_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1448_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1449_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1449_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_145_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_145_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1450_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1450_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1451_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1451_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1452_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1452_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1453_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1453_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1454_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1454_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1455_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1455_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1456_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1456_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1457_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1457_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1458_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1458_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1459_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1459_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_146_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_146_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1460_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1460_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1461_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1461_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1462_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1462_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1463_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1463_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1464_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1464_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1465_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1465_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1466_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1466_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1467_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1467_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1468_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1468_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1469_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1469_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_147_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_147_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1470_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1470_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1471_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1471_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1472_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1472_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1473_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1473_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1474_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1474_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1475_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1475_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1476_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1476_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1477_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1477_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1478_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1478_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1479_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1479_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_148_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_148_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1480_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1480_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1481_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1481_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1482_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1482_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1483_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1483_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1484_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1484_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1485_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1485_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1486_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1486_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1487_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2570 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1487_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1488_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1488_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1489_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1489_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_149_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_149_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1490_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1490_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1491_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1491_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1492_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1492_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1493_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1493_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1494_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1494_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1495_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1495_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1496_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1496_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1497_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1497_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1498_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1498_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1499_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1499_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_15_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_15_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_150_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_150_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1500_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1500_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1501_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1501_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1502_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1502_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1503_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2589 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1503_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1504_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1504_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1505_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1505_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1506_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1506_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1507_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1507_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1508_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1508_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1509_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1509_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_151_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_151_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1510_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1510_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1511_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1511_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1512_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1512_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1513_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1513_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1514_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1514_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1515_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1515_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1516_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1516_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1517_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1517_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1518_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1518_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1519_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2609 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1519_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_152_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_152_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1520_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1520_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1521_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1521_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1522_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1522_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1523_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1523_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1524_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1524_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1525_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1525_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1526_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1526_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1527_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1527_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1528_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1528_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1529_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1529_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_153_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_153_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1530_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1530_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1531_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1531_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1532_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1532_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1533_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1533_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1534_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1534_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1535_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2627 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1535_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1536_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_2718 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1536_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1537_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1537_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1538_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1538_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1539_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1539_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_154_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_154_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1540_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1540_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1541_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1541_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1542_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1542_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1543_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1543_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1544_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1544_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1545_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1545_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1546_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1546_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1547_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1547_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1548_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1548_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1549_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1549_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_155_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_155_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1550_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1550_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1551_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1551_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1552_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1552_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1553_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1553_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1554_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1554_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1555_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1555_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1556_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1556_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1557_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1557_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1558_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1558_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1559_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1559_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_156_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_156_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1560_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1560_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1561_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1561_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1562_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1562_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1563_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1563_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1564_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1564_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1565_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1565_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1566_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1566_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1567_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1567_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1568_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1568_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1569_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1569_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_157_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_157_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1570_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1570_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1571_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1571_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1572_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1572_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1573_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1573_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1574_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1574_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1575_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1575_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1576_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1576_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1577_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1577_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1578_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1578_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1579_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1579_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_158_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_158_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1580_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1580_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1581_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1581_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1582_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1582_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1583_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1583_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1584_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1584_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1585_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1585_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1586_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1586_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1587_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1587_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1588_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1588_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1589_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1589_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_159_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_159_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1590_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1590_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1591_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1591_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1592_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1592_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1593_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1593_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1594_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1594_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1595_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1595_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1596_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1596_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1597_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1597_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1598_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1598_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1599_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1599_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_16_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_16_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_160_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_160_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1600_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1600_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1601_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1601_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1602_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1602_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1603_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1603_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1604_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1604_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1605_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1605_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1606_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1606_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1607_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1607_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1608_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1608_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1609_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1609_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_161_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_161_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1610_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1610_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1611_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1611_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1612_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1612_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1613_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1613_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1614_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1614_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1615_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2718 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1615_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1616_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1616_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1617_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1617_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1618_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1618_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1619_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1619_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_162_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_162_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1620_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1620_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1621_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1621_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1622_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1622_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1623_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1623_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1624_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1624_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1625_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1625_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1626_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1626_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1627_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1627_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1628_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1628_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1629_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1629_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_163_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_163_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1630_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1630_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1631_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2738 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1631_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1632_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1632_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1633_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1633_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1634_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1634_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1635_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1635_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1636_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1636_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1637_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1637_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1638_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1638_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1639_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1639_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_164_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_164_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1640_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1640_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1641_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1641_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1642_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1642_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1643_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1643_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1644_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1644_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1645_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1645_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1646_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1646_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1647_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2756 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1647_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1648_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1648_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1649_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1649_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_165_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_165_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1650_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1650_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1651_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1651_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1652_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1652_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1653_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1653_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1654_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1654_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1655_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1655_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1656_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1656_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1657_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1657_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1658_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1658_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1659_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1659_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_166_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_166_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1660_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1660_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1661_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1661_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1662_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1662_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1663_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2775 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1663_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1664_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_2867 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1664_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1665_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1665_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1666_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1666_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1667_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1667_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1668_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1668_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1669_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1669_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_167_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_167_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1670_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1670_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1671_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1671_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1672_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1672_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1673_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1673_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1674_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1674_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1675_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1675_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1676_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1676_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1677_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1677_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1678_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1678_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1679_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1679_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_168_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_168_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1680_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1680_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1681_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1681_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1682_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1682_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1683_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1683_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1684_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1684_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1685_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1685_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1686_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1686_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1687_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1687_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1688_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1688_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1689_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1689_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_169_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_169_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1690_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1690_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1691_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1691_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1692_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1692_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1693_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1693_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1694_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1694_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1695_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1695_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1696_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1696_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1697_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1697_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1698_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1698_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1699_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1699_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_17_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_17_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_170_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_170_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1700_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1700_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1701_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1701_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1702_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1702_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1703_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1703_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1704_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1704_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1705_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1705_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1706_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1706_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1707_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1707_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1708_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1708_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1709_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1709_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_171_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_171_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1710_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1710_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1711_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1711_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1712_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1712_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1713_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1713_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1714_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1714_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1715_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1715_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1716_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1716_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1717_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1717_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1718_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1718_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1719_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1719_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_172_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_172_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1720_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1720_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1721_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1721_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1722_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1722_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1723_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1723_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1724_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1724_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1725_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1725_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1726_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1726_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1727_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1727_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1728_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1728_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1729_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1729_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_173_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_173_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1730_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1730_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1731_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1731_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1732_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1732_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1733_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1733_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1734_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1734_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1735_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1735_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1736_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1736_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1737_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1737_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1738_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1738_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1739_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1739_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_174_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_174_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1740_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1740_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1741_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1741_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1742_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1742_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1743_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2867 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1743_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1744_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1744_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1745_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1745_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1746_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1746_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1747_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1747_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1748_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1748_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1749_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1749_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_175_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_175_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1750_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1750_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1751_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1751_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1752_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1752_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1753_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1753_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1754_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1754_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1755_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1755_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1756_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1756_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1757_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1757_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1758_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1758_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1759_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2886 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1759_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_176_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_176_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1760_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1760_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1761_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1761_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1762_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1762_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1763_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1763_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1764_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1764_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1765_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1765_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1766_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1766_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1767_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1767_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1768_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1768_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1769_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1769_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_177_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_177_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1770_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1770_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1771_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1771_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1772_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1772_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1773_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1773_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1774_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1774_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1775_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2904 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1775_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1776_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1776_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1777_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1777_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1778_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1778_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1779_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1779_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_178_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_178_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1780_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1780_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1781_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1781_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1782_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1782_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1783_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1783_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1784_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1784_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1785_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1785_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1786_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1786_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1787_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1787_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1788_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1788_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1789_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1789_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_179_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_179_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1790_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1790_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1791_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2924 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_1791_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_18_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_18_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_180_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_180_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_181_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_181_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_182_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_182_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_183_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_183_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_184_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_184_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_185_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_185_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_186_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_186_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_187_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_187_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_188_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_188_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_189_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_189_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_19_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_19_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_190_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_190_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_191_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_191_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_192_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_192_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_193_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_193_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_194_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_194_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_195_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_195_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_196_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_196_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_197_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_197_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_198_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_198_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_199_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_199_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_2_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_2_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_20_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_20_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_200_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_200_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_201_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_201_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_202_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_202_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_203_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_203_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_204_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_204_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_205_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_205_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_206_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_206_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_207_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2419 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_207_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_208_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_208_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_209_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_209_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_21_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_21_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_210_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_210_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_211_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_211_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_212_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_212_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_213_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_213_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_214_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_214_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_215_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_215_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_216_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_216_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_217_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_217_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_218_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_218_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_219_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_219_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_22_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_22_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_220_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_220_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_221_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_221_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_222_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_222_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_223_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2607 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_223_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_224_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_224_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_225_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_225_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_226_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_226_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_227_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_227_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_228_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_228_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_229_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_229_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_23_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_23_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_230_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_230_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_231_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_231_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_232_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_232_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_233_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_233_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_234_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_234_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_235_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_235_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_236_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_236_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_237_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_237_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_238_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_238_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_239_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2795 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_239_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_24_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_24_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_240_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_240_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_241_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_241_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_242_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_242_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_243_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_243_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_244_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_244_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_245_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_245_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_246_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_246_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_247_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_247_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_248_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_248_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_249_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_249_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_25_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_25_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_250_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_250_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_251_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_251_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_252_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_252_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_253_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_253_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_254_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_254_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_255_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2977 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_255_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_256_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_3100 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_256_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_257_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_257_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_258_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_258_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_259_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_259_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_26_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_26_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_260_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_260_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_261_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_261_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_262_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_262_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_263_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_263_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_264_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_264_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_265_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_265_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_266_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_266_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_267_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_267_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_268_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_268_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_269_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_269_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_27_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_27_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_270_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_270_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_271_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_271_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_272_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_272_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_273_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_273_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_274_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_274_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_275_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_275_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_276_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_276_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_277_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_277_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_278_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_278_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_279_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_279_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_28_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_28_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_280_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_280_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_281_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_281_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_282_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_282_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_283_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_283_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_284_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_284_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_285_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_285_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_286_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_286_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_287_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_287_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_288_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_288_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_289_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_289_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_29_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_29_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_290_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_290_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_291_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_291_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_292_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_292_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_293_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_293_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_294_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_294_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_295_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_295_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_296_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_296_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_297_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_297_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_298_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_298_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_299_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_299_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_3_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_3_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_30_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_30_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_300_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_300_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_301_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_301_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_302_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_302_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_303_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_303_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_304_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_304_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_305_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_305_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_306_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_306_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_307_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_307_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_308_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_308_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_309_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_309_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_31_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_31_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_310_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_310_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_311_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_311_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_312_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_312_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_313_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_313_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_314_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_314_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_315_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_315_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_316_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_316_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_317_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_317_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_318_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_318_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_319_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_319_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_32_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_32_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_320_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_320_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_321_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_321_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_322_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_322_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_323_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_323_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_324_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_324_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_325_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_325_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_326_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_326_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_327_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_327_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_328_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_328_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_329_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_329_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_33_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_33_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_330_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_330_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_331_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_331_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_332_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_332_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_333_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_333_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_334_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_334_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_335_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3100 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_335_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_336_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_336_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_337_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_337_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_338_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_338_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_339_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_339_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_34_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_34_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_340_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_340_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_341_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_341_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_342_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_342_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_343_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_343_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_344_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_344_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_345_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_345_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_346_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_346_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_347_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_347_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_348_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_348_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_349_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_349_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_35_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_35_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_350_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_350_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_351_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3119 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_351_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_352_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_352_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_353_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_353_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_354_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_354_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_355_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_355_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_356_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_356_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_357_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_357_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_358_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_358_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_359_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_359_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_36_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_36_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_360_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_360_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_361_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_361_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_362_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_362_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_363_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_363_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_364_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_364_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_365_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_365_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_366_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_366_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_367_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3137 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_367_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_368_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_368_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_369_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_369_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_37_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_37_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_370_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_370_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_371_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_371_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_372_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_372_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_373_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_373_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_374_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_374_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_375_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_375_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_376_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_376_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_377_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_377_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_378_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_378_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_379_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_379_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_38_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_38_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_380_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_380_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_381_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_381_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_382_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_382_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_383_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3157 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_383_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_384_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_3246 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_384_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_385_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_385_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_386_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_386_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_387_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_387_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_388_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_388_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_389_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_389_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_39_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_39_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_390_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_390_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_391_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_391_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_392_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_392_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_393_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_393_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_394_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_394_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_395_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_395_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_396_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_396_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_397_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_397_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_398_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_398_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_399_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_399_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_4_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_4_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_40_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_40_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_400_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_400_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_401_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_401_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_402_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_402_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_403_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_403_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_404_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_404_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_405_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_405_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_406_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_406_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_407_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_407_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_408_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_408_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_409_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_409_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_41_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_41_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_410_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_410_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_411_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_411_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_412_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_412_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_413_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_413_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_414_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_414_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_415_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_415_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_416_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_416_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_417_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_417_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_418_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_418_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_419_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_419_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_42_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_42_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_420_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_420_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_421_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_421_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_422_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_422_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_423_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_423_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_424_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_424_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_425_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_425_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_426_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_426_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_427_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_427_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_428_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_428_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_429_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_429_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_43_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_43_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_430_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_430_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_431_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_431_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_432_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_432_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_433_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_433_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_434_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_434_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_435_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_435_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_436_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_436_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_437_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_437_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_438_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_438_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_439_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_439_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_44_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_44_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_440_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_440_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_441_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_441_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_442_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_442_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_443_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_443_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_444_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_444_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_445_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_445_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_446_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_446_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_447_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_447_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_448_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_448_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_449_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_449_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_45_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_45_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_450_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_450_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_451_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_451_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_452_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_452_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_453_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_453_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_454_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_454_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_455_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_455_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_456_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_456_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_457_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_457_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_458_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_458_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_459_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_459_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_46_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_46_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_460_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_460_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_461_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_461_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_462_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_462_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_463_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3246 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_463_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_464_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_464_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_465_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_465_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_466_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_466_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_467_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_467_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_468_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_468_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_469_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_469_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_47_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_47_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_470_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_470_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_471_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_471_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_472_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_472_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_473_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_473_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_474_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_474_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_475_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_475_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_476_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_476_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_477_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_477_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_478_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_478_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_479_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3266 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_479_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_48_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_48_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_480_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_480_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_481_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_481_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_482_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_482_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_483_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_483_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_484_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_484_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_485_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_485_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_486_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_486_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_487_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_487_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_488_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_488_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_489_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_489_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_49_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_49_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_490_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_490_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_491_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_491_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_492_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_492_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_493_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_493_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_494_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_494_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_495_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3284 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_495_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_496_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_496_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_497_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_497_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_498_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_498_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_499_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_499_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_5_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_5_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_50_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_50_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_500_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_500_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_501_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_501_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_502_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_502_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_503_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_503_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_504_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_504_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_505_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_505_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_506_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_506_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_507_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_507_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_508_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_508_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_509_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_509_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_51_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_51_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_510_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_510_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_511_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3303 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_511_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_512_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_3393 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_512_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_513_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_513_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_514_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_514_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_515_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_515_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_516_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_516_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_517_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_517_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_518_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_518_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_519_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_519_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_52_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_52_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_520_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_520_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_521_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_521_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_522_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_522_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_523_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_523_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_524_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_524_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_525_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_525_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_526_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_526_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_527_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_527_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_528_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_528_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_529_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_529_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_53_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_53_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_530_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_530_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_531_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_531_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_532_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_532_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_533_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_533_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_534_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_534_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_535_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_535_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_536_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_536_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_537_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_537_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_538_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_538_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_539_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_539_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_54_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_54_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_540_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_540_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_541_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_541_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_542_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_542_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_543_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_543_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_544_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_544_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_545_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_545_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_546_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_546_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_547_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_547_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_548_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_548_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_549_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_549_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_55_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_55_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_550_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_550_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_551_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_551_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_552_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_552_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_553_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_553_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_554_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_554_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_555_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_555_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_556_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_556_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_557_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_557_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_558_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_558_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_559_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_559_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_56_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_56_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_560_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_560_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_561_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_561_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_562_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_562_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_563_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_563_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_564_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_564_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_565_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_565_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_566_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_566_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_567_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_567_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_568_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_568_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_569_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_569_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_57_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_57_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_570_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_570_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_571_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_571_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_572_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_572_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_573_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_573_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_574_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_574_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_575_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_575_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_576_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_576_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_577_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_577_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_578_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_578_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_579_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_579_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_58_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_58_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_580_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_580_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_581_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_581_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_582_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_582_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_583_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_583_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_584_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_584_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_585_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_585_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_586_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_586_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_587_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_587_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_588_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_588_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_589_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_589_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_59_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_59_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_590_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_590_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_591_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3393 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_591_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_592_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_592_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_593_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_593_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_594_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_594_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_595_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_595_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_596_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_596_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_597_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_597_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_598_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_598_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_599_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_599_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_6_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_6_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_60_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_60_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_600_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_600_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_601_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_601_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_602_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_602_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_603_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_603_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_604_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_604_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_605_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_605_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_606_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_606_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_607_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3411 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_607_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_608_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_608_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_609_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_609_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_61_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_61_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_610_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_610_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_611_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_611_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_612_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_612_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_613_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_613_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_614_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_614_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_615_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_615_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_616_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_616_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_617_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_617_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_618_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_618_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_619_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_619_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_62_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_62_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_620_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_620_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_621_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_621_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_622_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_622_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_623_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3430 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_623_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_624_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_624_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_625_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_625_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_626_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_626_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_627_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_627_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_628_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_628_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_629_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_629_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_63_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2234 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_63_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_630_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_630_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_631_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_631_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_632_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_632_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_633_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_633_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_634_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_634_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_635_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_635_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_636_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_636_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_637_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_637_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_638_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_638_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_639_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3449 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_639_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_64_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_64_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_640_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_3539 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_640_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_641_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_641_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_642_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_642_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_643_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_643_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_644_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_644_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_645_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_645_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_646_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_646_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_647_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_647_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_648_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_648_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_649_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_649_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_65_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_65_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_650_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_650_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_651_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_651_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_652_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_652_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_653_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_653_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_654_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_654_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_655_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_655_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_656_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_656_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_657_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_657_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_658_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_658_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_659_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_659_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_66_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_66_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_660_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_660_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_661_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_661_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_662_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_662_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_663_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_663_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_664_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_664_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_665_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_665_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_666_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_666_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_667_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_667_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_668_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_668_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_669_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_669_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_67_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_67_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_670_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_670_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_671_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_671_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_672_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_672_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_673_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_673_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_674_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_674_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_675_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_675_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_676_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_676_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_677_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_677_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_678_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_678_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_679_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_679_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_68_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_68_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_680_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_680_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_681_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_681_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_682_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_682_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_683_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_683_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_684_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_684_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_685_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_685_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_686_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_686_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_687_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_687_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_688_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_688_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_689_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_689_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_69_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_69_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_690_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_690_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_691_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_691_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_692_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_692_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_693_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_693_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_694_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_694_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_695_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_695_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_696_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_696_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_697_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_697_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_698_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_698_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_699_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_699_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_7_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_7_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_70_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_70_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_700_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_700_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_701_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_701_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_702_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_702_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_703_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_703_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_704_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_704_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_705_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_705_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_706_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_706_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_707_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_707_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_708_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_708_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_709_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_709_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_71_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_71_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_710_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_710_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_711_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_711_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_712_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_712_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_713_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_713_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_714_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_714_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_715_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_715_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_716_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_716_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_717_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_717_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_718_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_718_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_719_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3539 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_719_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_72_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_72_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_720_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_720_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_721_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_721_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_722_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_722_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_723_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_723_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_724_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_724_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_725_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_725_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_726_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_726_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_727_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_727_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_728_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_728_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_729_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_729_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_73_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_73_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_730_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_730_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_731_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_731_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_732_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_732_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_733_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_733_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_734_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_734_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_735_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3557 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_735_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_736_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_736_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_737_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_737_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_738_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_738_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_739_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_739_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_74_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_74_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_740_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_740_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_741_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_741_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_742_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_742_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_743_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_743_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_744_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_744_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_745_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_745_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_746_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_746_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_747_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_747_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_748_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_748_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_749_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_749_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_75_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_75_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_750_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_750_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_751_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3576 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_751_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_752_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_752_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_753_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_753_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_754_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_754_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_755_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_755_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_756_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_756_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_757_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_757_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_758_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_758_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_759_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_759_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_76_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_76_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_760_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_760_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_761_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_761_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_762_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_762_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_763_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_763_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_764_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_764_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_765_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_765_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_766_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_766_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_767_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3594 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_767_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_768_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_3684 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_768_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_769_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_769_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_77_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_77_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_770_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_770_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_771_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_771_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_772_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_772_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_773_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_773_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_774_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_774_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_775_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_775_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_776_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_776_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_777_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_777_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_778_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_778_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_779_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_779_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_78_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_78_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_780_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_780_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_781_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_781_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_782_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_782_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_783_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_783_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_784_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_784_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_785_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_785_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_786_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_786_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_787_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_787_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_788_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_788_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_789_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_789_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_79_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_79_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_790_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_790_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_791_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_791_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_792_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_792_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_793_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_793_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_794_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_794_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_795_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_795_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_796_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_796_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_797_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_797_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_798_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_798_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_799_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_799_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_8_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_8_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_80_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_80_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_800_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_800_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_801_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_801_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_802_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_802_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_803_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_803_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_804_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_804_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_805_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_805_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_806_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_806_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_807_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_807_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_808_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_808_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_809_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_809_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_81_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_81_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_810_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_810_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_811_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_811_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_812_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_812_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_813_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_813_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_814_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_814_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_815_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_815_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_816_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_816_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_817_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_817_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_818_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_818_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_819_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_819_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_82_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_82_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_820_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_820_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_821_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_821_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_822_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_822_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_823_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_823_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_824_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_824_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_825_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_825_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_826_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_826_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_827_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_827_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_828_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_828_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_829_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_829_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_83_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_83_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_830_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_830_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_831_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_831_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_832_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_832_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_833_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_833_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_834_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_834_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_835_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_835_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_836_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_836_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_837_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_837_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_838_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_838_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_839_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_839_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_84_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_84_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_840_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_840_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_841_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_841_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_842_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_842_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_843_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_843_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_844_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_844_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_845_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_845_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_846_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_846_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_847_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3684 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_847_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_848_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_848_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_849_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_849_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_85_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_85_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_850_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_850_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_851_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_851_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_852_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_852_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_853_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_853_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_854_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_854_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_855_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_855_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_856_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_856_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_857_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_857_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_858_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_858_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_859_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_859_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_86_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_86_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_860_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_860_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_861_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_861_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_862_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_862_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_863_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3703 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_863_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_864_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_864_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_865_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_865_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_866_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_866_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_867_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_867_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_868_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_868_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_869_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_869_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_87_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_87_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_870_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_870_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_871_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_871_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_872_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_872_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_873_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_873_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_874_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_874_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_875_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_875_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_876_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_876_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_877_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_877_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_878_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_878_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_879_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3723 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_879_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_88_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_88_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_880_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_880_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_881_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_881_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_882_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_882_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_883_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_883_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_884_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_884_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_885_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_885_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_886_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_886_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_887_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_887_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_888_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_888_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_889_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_889_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_89_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_89_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_890_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_890_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_891_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_891_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_892_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_892_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_893_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_893_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_894_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_894_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_895_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3741 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_895_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_896_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (~(or_dcpl_3830 | or_dcpl_2030)) & (fsm_output[2]) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_896_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_897_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_897_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_898_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_898_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_899_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_899_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_9_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2035 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_9_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_90_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_90_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_900_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_900_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_901_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_901_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_902_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_902_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_903_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_903_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_904_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_904_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_905_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_905_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_906_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_906_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_907_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_907_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_908_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_908_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_909_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_909_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_91_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_91_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_910_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_910_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_911_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_911_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_912_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_912_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_913_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_913_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_914_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_914_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_915_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_915_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_916_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_916_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_917_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_917_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_918_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_918_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_919_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_919_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_92_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_92_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_920_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_920_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_921_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_921_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_922_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_922_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_923_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_923_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_924_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_924_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_925_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_925_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_926_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_926_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_927_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_927_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_928_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_928_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_929_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_929_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_93_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_93_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_930_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_930_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_931_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_931_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_932_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_932_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_933_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_933_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_934_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_934_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_935_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_935_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_936_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_936_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_937_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_937_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_938_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_938_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_939_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_939_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_94_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_94_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_940_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_940_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_941_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_941_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_942_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_942_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_943_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_943_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_944_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2030)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_944_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_945_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2038)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_945_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_946_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2110)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_946_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_947_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2113)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_947_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_948_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2115)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_948_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_949_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2117)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_949_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_95_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2793 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_95_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_950_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2120)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_950_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_951_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2122)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_951_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_952_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2124)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_952_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_953_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2126)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_953_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_954_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2043)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_954_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_955_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2129)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_955_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_956_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2131)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_956_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_957_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2133)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_957_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_958_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2135)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_958_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_959_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2081 | or_dcpl_2137)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_959_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_96_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_96_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_960_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_960_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_961_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_961_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_962_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_962_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_963_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_963_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_964_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_964_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_965_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_965_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_966_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_966_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_967_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_967_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_968_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_968_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_969_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_969_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_97_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_97_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_970_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_970_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_971_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_971_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_972_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_972_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_973_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_973_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_974_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_974_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_975_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3830 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_975_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_976_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_976_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_977_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_977_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_978_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_978_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_979_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_979_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_98_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_98_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_980_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_980_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_981_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_981_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_982_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_982_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_983_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_983_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_984_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2052)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_984_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_985_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2060)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_985_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_986_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2064)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_986_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_987_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2067)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_987_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_988_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2070)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_988_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_989_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2072)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_989_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_99_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2050 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_99_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_990_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2074)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_990_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_991_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_3850 | or_dcpl_2076)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_991_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_992_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2078)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_992_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_993_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2083)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_993_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_994_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2087)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_994_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_995_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2089)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_995_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_996_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2048)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_996_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_997_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2085)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_997_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_998_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2093)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_998_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_999_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[2]) & (~(or_dcpl_2057 | or_dcpl_2095)) ) begin
      nnet_dense_latency_input_t_layer2_t_config2_mult_999_lpi_3 <= z_out_5_19_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_0_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[1]) | (fsm_output[3]) | and_5052_rgt | or_6921_rgt | and_5057_rgt
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_0_lpi_3 <= MUX1HOT_v_16_4_2(Product1_mux_nl,
          16'b0000001001000000, z_out_6, 16'b0000000010000000, {(fsm_output[1]) ,
          (fsm_output[3]) , nnet_dense_latency_input_t_layer2_t_config2_acc_or_nl
          , or_6921_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Result_ires_7_0_sva_1 <= 8'b00000000;
    end
    else if ( ~((fsm_output[14]) | (fsm_output[0]) | (fsm_output[13]) | (fsm_output[9]))
        ) begin
      Result_ires_7_0_sva_1 <= MUX_v_8_2_2(({1'b0 , mux_nl}), z_out_2, fsm_output[8]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_127_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_127_lpi_3 <= MUX_v_16_2_2(16'b1111110110000000,
          z_out_6, and_5067_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_126_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_126_lpi_3 <= MUX_v_16_2_2(16'b1111111001000000,
          z_out_6, and_5074_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_1_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[3]) | and_5081_rgt | or_tmp_2362 | and_5086_rgt ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_1_lpi_3 <= MUX1HOT_v_16_3_2(16'b0000001011000000,
          z_out_6, 16'b1111111100000000, {(fsm_output[3]) , nnet_dense_latency_input_t_layer2_t_config2_acc_or_4_nl
          , or_tmp_2362});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_125_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_125_lpi_3 <= MUX_v_16_2_2(16'b1111111001000000,
          z_out_6, and_5095_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_2_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4424 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_2_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5102_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_124_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_124_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5109_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_3_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4424 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_3_lpi_3 <= MUX_v_16_2_2(16'b1111110110000000,
          z_out_6, and_5116_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_123_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_123_lpi_3 <= MUX_v_16_2_2(16'b0000000101000000,
          z_out_6, and_5123_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_4_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4399 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_4_lpi_3 <= MUX_v_16_2_2(16'b0000000100000000,
          z_out_6, and_5130_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_122_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_122_lpi_3 <= MUX_v_16_2_2(16'b1111110010000000,
          z_out_6, and_5137_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_5_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4399 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_5_lpi_3 <= MUX_v_16_2_2(16'b1111111110000000,
          z_out_6, and_5144_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_121_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_121_lpi_3 <= MUX_v_16_2_2(16'b0000000110000000,
          z_out_6, and_5151_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_6_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4424 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_6_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5158_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_120_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_120_lpi_3 <= MUX_v_16_2_2(16'b0000000100000000,
          z_out_6, and_5165_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_7_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4424 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_7_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5172_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_119_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_119_lpi_3 <= MUX_v_16_2_2(16'b1111111110000000,
          z_out_6, and_5179_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_8_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4399 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_8_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5186_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_118_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_118_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5193_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_9_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4399 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_9_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5200_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_117_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_117_lpi_3 <= MUX_v_16_2_2(16'b0000000010000000,
          z_out_6, and_5207_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_10_lpi_3 <= 16'b0000000000000000;
    end
    else if ( (fsm_output[3]) | and_5214_rgt | or_tmp_2362 | and_5219_rgt ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_10_lpi_3 <= MUX1HOT_v_16_3_2(16'b0000000110000000,
          z_out_6, 16'b0000000011000000, {(fsm_output[3]) , nnet_dense_latency_input_t_layer2_t_config2_acc_or_23_nl
          , or_tmp_2362});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_116_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_116_lpi_3 <= MUX_v_16_2_2(16'b0000000011000000,
          z_out_6, and_5228_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_11_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4424 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_11_lpi_3 <= MUX_v_16_2_2(16'b1111111001000000,
          z_out_6, and_5235_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_115_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_115_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5242_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_12_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4399 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_12_lpi_3 <= MUX_v_16_2_2(16'b0000000100000000,
          z_out_6, and_5249_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_114_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4412 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_114_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5256_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_13_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4399 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_13_lpi_3 <= MUX_v_16_2_2(16'b1111111110000000,
          z_out_6, and_5263_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_113_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_113_lpi_3 <= MUX_v_16_2_2(16'b0000001101000000,
          z_out_6, and_5270_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_14_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4424 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_14_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5277_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_112_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4422 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_112_lpi_3 <= MUX_v_16_2_2(16'b0000000101000000,
          z_out_6, and_5284_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_15_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4424 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_15_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5291_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_111_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_111_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5298_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_16_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_16_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5305_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_110_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_110_lpi_3 <= nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_17_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_17_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5319_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_109_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_109_lpi_3 <= nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_18_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_18_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5333_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_108_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_108_lpi_3 <= MUX_v_16_2_2(16'b1111111001000000,
          z_out_6, and_5340_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_19_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_19_lpi_3 <= nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_107_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_107_lpi_3 <= MUX_v_16_2_2(16'b0000000100000000,
          z_out_6, and_5354_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_20_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_20_lpi_3 <= MUX_v_16_2_2(16'b1111111101000000,
          z_out_6, and_5361_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_106_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_106_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5368_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_21_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_21_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5375_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_105_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_105_lpi_3 <= MUX_v_16_2_2(16'b0000001010000000,
          z_out_6, and_5382_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_22_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_22_lpi_3 <= MUX_v_16_2_2(16'b0000000101000000,
          z_out_6, and_5389_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_104_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_104_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5396_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_23_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_23_lpi_3 <= MUX_v_16_2_2(16'b1111111101000000,
          z_out_6, and_5403_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_103_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_103_lpi_3 <= MUX_v_16_2_2(16'b1111111001000000,
          z_out_6, and_5410_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_24_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_24_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5417_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_102_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_102_lpi_3 <= MUX_v_16_2_2(16'b1111110110000000,
          z_out_6, and_5424_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_25_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_25_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5431_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_101_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_101_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5438_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_26_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_26_lpi_3 <= MUX_v_16_2_2(16'b0000001100000000,
          z_out_6, and_5445_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_100_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_100_lpi_3 <= MUX1HOT_v_16_3_2(16'b1111111110000000,
          z_out_6, layer6_out_rsci_idat_15_0, {(fsm_output[3]) , and_5452_nl , (fsm_output[14])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_27_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_27_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5461_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_99_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_99_lpi_3 <= MUX_v_16_2_2(16'b1111111110000000,
          z_out_6, and_5468_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_28_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_28_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5475_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_98_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4457 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_98_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5482_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_29_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4460 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_29_lpi_3 <= MUX_v_16_2_2(16'b1111110101000000,
          z_out_6, and_5489_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_97_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_97_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5496_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_30_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_30_lpi_3 <= MUX_v_16_2_2(16'b0000000011000000,
          z_out_6, and_5503_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_96_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4464 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_96_lpi_3 <= MUX_v_16_2_2(16'b0000000011000000,
          z_out_6, and_5510_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_31_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4466 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_31_lpi_3 <= MUX_v_16_2_2(16'b0000001100000000,
          z_out_6, and_5517_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_95_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_95_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5524_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_32_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_32_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5531_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_94_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_94_lpi_3 <= MUX_v_16_2_2(16'b0000001001000000,
          z_out_6, and_5538_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_33_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_33_lpi_3 <= MUX_v_16_2_2(16'b0000001001000000,
          z_out_6, and_5545_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_93_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_93_lpi_3 <= MUX_v_16_2_2(16'b0000000111000000,
          z_out_6, and_5552_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_34_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_34_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5559_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_92_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_92_lpi_3 <= MUX_v_16_2_2(16'b1111111001000000,
          z_out_6, and_5566_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_35_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_35_lpi_3 <= nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_91_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_91_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5580_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_36_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_36_lpi_3 <= MUX_v_16_2_2(16'b0000000010000000,
          z_out_6, and_5587_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_90_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_90_lpi_3 <= MUX_v_16_2_2(16'b1111111101000000,
          z_out_6, and_5594_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_37_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_37_lpi_3 <= MUX_v_16_2_2(16'b0000001000000000,
          z_out_6, and_5601_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_89_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_89_lpi_3 <= MUX_v_16_2_2(16'b1111111101000000,
          z_out_6, and_5608_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_38_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_38_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5615_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_88_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_88_lpi_3 <= nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_39_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_39_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5629_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_87_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_87_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5636_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_40_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_40_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5643_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_86_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_86_lpi_3 <= MUX_v_16_2_2(16'b0000000100000000,
          z_out_6, and_5650_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_41_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_41_lpi_3 <= MUX_v_16_2_2(16'b0000001000000000,
          z_out_6, and_5657_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_85_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_85_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5664_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_42_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_42_lpi_3 <= MUX_v_16_2_2(16'b1111111101000000,
          z_out_6, and_5671_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_84_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_84_lpi_3 <= MUX_v_16_2_2(16'b1111111110000000,
          z_out_6, and_5678_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_43_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_43_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5685_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_83_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_83_lpi_3 <= MUX_v_16_2_2(16'b0000001001000000,
          z_out_6, and_5692_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_44_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_44_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5699_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_82_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4494 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_82_lpi_3 <= MUX_v_16_2_2(16'b1111110110000000,
          z_out_6, and_5706_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_45_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4496 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_45_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5713_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_81_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_81_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5720_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_46_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_46_lpi_3 <= MUX_v_16_2_2(16'b1111111110000000,
          z_out_6, and_5727_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_80_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4500 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_80_lpi_3 <= MUX_v_16_2_2(16'b0000000011000000,
          z_out_6, and_5734_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_47_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4502 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_47_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5741_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_79_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_79_lpi_3 <= MUX_v_16_2_2(16'b0000000011000000,
          z_out_6, and_5748_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_48_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_48_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5755_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_78_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_78_lpi_3 <= nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_49_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_49_lpi_3 <= MUX_v_16_2_2(16'b0000000110000000,
          z_out_6, and_5769_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_77_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_77_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5776_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_50_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_50_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5783_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_76_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_76_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5790_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_51_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_51_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5797_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_75_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_75_lpi_3 <= MUX_v_16_2_2(16'b1111111110000000,
          z_out_6, and_5804_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_52_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_52_lpi_3 <= MUX_v_16_2_2(16'b0000001000000000,
          z_out_6, and_5811_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_74_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_74_lpi_3 <= MUX_v_16_2_2(16'b1111110111000000,
          z_out_6, and_5818_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_53_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_53_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5825_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_73_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_73_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5832_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_54_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_54_lpi_3 <= MUX_v_16_2_2(16'b0000001001000000,
          z_out_6, and_5839_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_72_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_72_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5846_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_55_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_55_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5853_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_71_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_71_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5860_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_56_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_56_lpi_3 <= MUX_v_16_2_2(16'b1111111000000000,
          z_out_6, and_5867_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_70_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_70_lpi_3 <= MUX_v_16_2_2(16'b0000000111000000,
          z_out_6, and_5874_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_57_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_57_lpi_3 <= MUX_v_16_2_2(16'b0000000100000000,
          z_out_6, and_5881_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_69_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4434) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_69_lpi_3 <= MUX_v_16_2_2(16'b0000000011000000,
          z_out_6, and_5888_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_58_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4432) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_58_lpi_3 <= MUX_v_16_2_2(16'b1111110110000000,
          z_out_6, and_5895_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_68_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4430) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_68_lpi_3 <= MUX_v_16_2_2(16'b1111111111000000,
          z_out_6, and_5902_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_59_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4428) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_59_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5909_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_67_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_67_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5916_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_60_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_60_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5923_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_66_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4530 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_66_lpi_3 <= MUX_v_16_2_2(16'b1111111011000000,
          z_out_6, and_5930_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_61_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4532 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_61_lpi_3 <= MUX_v_16_2_2(16'b0000000001000000,
          z_out_6, and_5937_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_65_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4420) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_65_lpi_3 <= MUX_v_16_2_2(16'b1111111010000000,
          z_out_6, and_5944_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_62_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4415) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_62_lpi_3 <= MUX_v_16_2_2(16'b1111111100000000,
          z_out_6, and_5951_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_64_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4536 | or_dcpl_4397) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_64_lpi_3 <= MUX_v_16_2_2(16'b1111110010000000,
          z_out_6, and_5958_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_63_lpi_3 <= 16'b0000000000000000;
    end
    else if ( ~(and_5068_cse | ((or_dcpl_4538 | or_dcpl_4410) & (fsm_output[4])))
        ) begin
      nnet_dense_latency_input_t_layer2_t_config2_acc_63_lpi_3 <= nnet_dense_latency_input_t_layer2_t_config2_acc_nnet_dense_latency_input_t_layer2_t_config2_acc_and_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Product1_1_ii_7_0_sva_6_0 <= 7'b0000000;
    end
    else if ( Product1_1_ii_or_cse ) begin
      Product1_1_ii_7_0_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (z_out_2[6:0]), (fsm_output[10]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1 <= 8'b00000000;
    end
    else if ( nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_or_cse | (fsm_output[7])
        | nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1_mx0c2 ) begin
      nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1 <= MUX1HOT_v_8_3_2(({1'b0
          , and_nl}), z_out_2, ({6'b000000 , Product2_1_jj_Product2_1_jj_and_1_nl}),
          {nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_or_cse , (fsm_output[7])
          , nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1_mx0c2});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_7_0_sva_1 <= 8'b00000000;
    end
    else if ( nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_or_cse ) begin
      nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_7_0_sva_1 <= MUX_v_8_2_2(({1'b0
          , Product2_jj_Product2_jj_and_1_nl}), z_out_2, fsm_output[6]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer4_out_9_lpi_2_dfm <= 1'b0;
    end
    else if ( ~ or_tmp_2754 ) begin
      layer4_out_9_lpi_2_dfm <= ((Accum2_mux_131[9]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1)
          & operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer4_out_8_1_lpi_2_dfm <= 8'b00000000;
    end
    else if ( ~ or_tmp_2754 ) begin
      layer4_out_8_1_lpi_2_dfm <= MUX_v_8_2_2(8'b00000000, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl,
          operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer4_out_0_lpi_2_dfm <= 1'b0;
    end
    else if ( ~ or_tmp_2754 ) begin
      layer4_out_0_lpi_2_dfm <= ((Accum2_mux_131[0]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1)
          & operator_16_6_true_AC_RND_CONV_AC_SAT_acc_itm_16_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      Result_1_Result_1_nor_itm <= 1'b0;
    end
    else begin
      Result_1_Result_1_nor_itm <= ~((z_out_2[2]) | ((z_out_1[0]) ^ (z_out_1[1])));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_0_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_0_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_1_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_1_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_2_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_2_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_3_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_3_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_4_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_4_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_5_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_5_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_6_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_6_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_7_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_7_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_8_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_8_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_9_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_9_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_10_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_10_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_11_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_11_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_12_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_12_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_13_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_13_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_14_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_14_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_15_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_15_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_16_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_16_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_17_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_17_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_18_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_18_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_19_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_19_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_20_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_20_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_21_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_21_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_22_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_22_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_23_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_23_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_24_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_24_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_25_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_25_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_26_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_26_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_27_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_27_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_28_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_28_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_29_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_29_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_30_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_30_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_31_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_31_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_32_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_32_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_33_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_33_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_34_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_34_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_35_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_35_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_36_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_36_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_37_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_37_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_38_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_38_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_39_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_39_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_40_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_40_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_41_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_41_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_42_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_42_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_43_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_43_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_44_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_44_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_45_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_45_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_46_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_46_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_47_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_47_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_48_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_48_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_49_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_49_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_50_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_50_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_51_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_51_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_52_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_52_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_53_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_53_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_54_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_54_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_55_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_55_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_56_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_56_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_57_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_57_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_58_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_58_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_59_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_59_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_60_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_60_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_61_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_61_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_62_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_62_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_63_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_63_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_64_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_64_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_65_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_65_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_66_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_66_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_67_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_67_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_68_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_68_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_69_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_69_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_70_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_70_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_71_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_71_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_72_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_72_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_73_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_73_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_74_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_74_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_75_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_75_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_76_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_76_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_77_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_77_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_78_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_78_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_79_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_79_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_80_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_80_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_81_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_81_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_82_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_82_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_83_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_83_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_84_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_84_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_85_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_85_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_86_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_86_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_87_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_87_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_88_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_88_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_89_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_89_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_90_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_90_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_91_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_91_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_92_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_92_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_93_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_93_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_94_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_94_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_95_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_95_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_96_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_96_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_97_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_97_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_98_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_98_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_99_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_99_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_100_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_100_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_101_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_101_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_102_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_102_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_103_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_103_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_104_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_104_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_105_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_105_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_106_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_106_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_107_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_107_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_108_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_108_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_109_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_109_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_110_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_110_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_111_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_111_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_112_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_112_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_113_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3953 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_113_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_114_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_114_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_115_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3992 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_115_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_116_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_116_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_117_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3966 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_117_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_118_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_118_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_119_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3971 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_119_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_120_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_120_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_121_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3974 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_121_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_122_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_122_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_123_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3960 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_123_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_124_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_124_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_125_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3980 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_125_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_126_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_126_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_127_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_3984 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_127_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_128_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_128_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_129_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_129_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_130_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_130_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_131_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_131_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_132_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_132_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_133_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_133_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_134_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_134_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_135_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_135_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_136_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_136_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_137_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_137_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_138_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_138_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_139_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_139_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_140_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_140_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_141_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_141_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_142_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_142_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_143_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_143_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_144_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_144_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_145_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_145_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_146_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_146_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_147_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_147_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_148_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_148_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_149_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_149_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_150_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_150_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_151_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_151_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_152_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_152_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_153_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_153_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_154_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_154_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_155_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_155_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_156_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_156_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_157_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_157_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_158_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_158_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_159_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_159_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_160_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_160_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_161_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_161_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_162_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_162_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_163_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_163_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_164_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_164_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_165_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_165_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_166_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_166_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_167_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_167_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_168_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_168_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_169_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_169_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_170_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_170_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_171_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_171_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_172_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_172_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_173_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_173_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_174_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_174_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_175_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_175_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_176_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_176_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_177_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_177_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_178_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_178_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_179_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_179_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_180_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_180_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_181_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_181_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_182_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_182_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_183_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_183_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_184_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_184_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_185_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_185_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_186_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_186_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_187_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_187_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_188_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_188_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_189_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_189_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_190_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_190_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_191_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_191_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_192_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_192_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_193_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_193_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_194_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_194_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_195_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_195_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_196_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_196_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_197_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_197_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_198_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_198_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_199_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_199_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_200_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_200_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_201_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_201_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_202_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_202_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_203_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_203_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_204_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_204_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_205_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_205_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_206_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_206_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_207_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_207_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_208_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_208_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_209_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_209_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_210_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_210_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_211_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_211_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_212_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_212_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_213_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_213_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_214_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_214_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_215_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_215_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_216_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_216_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_217_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_217_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_218_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_218_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_219_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_219_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_220_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_220_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_221_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_221_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_222_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_222_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_223_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_223_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_224_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_224_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_225_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_225_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_226_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_226_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_227_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_227_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_228_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_228_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_229_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_229_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_230_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_230_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_231_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_231_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_232_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_232_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_233_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_233_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_234_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_234_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_235_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_235_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_236_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_236_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_237_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_237_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_238_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_238_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_239_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_239_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_240_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_240_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_241_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4010 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_241_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_242_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_242_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_243_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4015 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_243_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_244_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_244_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_245_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4018 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_245_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_246_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_246_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_247_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4021 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_247_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_248_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_248_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_249_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4024 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_249_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_250_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_250_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_251_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4027 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_251_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_252_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_252_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_253_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4031 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_253_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_254_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_254_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_255_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4034 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_255_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_256_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_256_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_257_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_257_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_258_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_258_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_259_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_259_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_260_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_260_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_261_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_261_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_262_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_262_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_263_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_263_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_264_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_264_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_265_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_265_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_266_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_266_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_267_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_267_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_268_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_268_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_269_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_269_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_270_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_3949) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_270_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_271_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_3956) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_271_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_272_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_272_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_273_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_273_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_274_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_274_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_275_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_275_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_276_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_276_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_277_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_277_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_278_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_278_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_279_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_279_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_280_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_280_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_281_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_281_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_282_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_282_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_283_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_283_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_284_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_284_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_285_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_285_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_286_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4038) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_286_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_287_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4040) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_287_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_288_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_288_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_289_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_289_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_290_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_290_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_291_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_291_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_292_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_292_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_293_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_293_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_294_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_294_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_295_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_295_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_296_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_296_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_297_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_297_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_298_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_298_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_299_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_299_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_300_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_300_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_301_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_301_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_302_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4058) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_302_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_303_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4060) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_303_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_304_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_304_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_305_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_305_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_306_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_306_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_307_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_307_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_308_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_308_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_309_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_309_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_310_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_310_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_311_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_311_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_312_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_312_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_313_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_313_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_314_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_314_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_315_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_315_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_316_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_316_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_317_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_317_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_318_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4077) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_318_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_319_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4079) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_319_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_320_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_320_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_321_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_321_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_322_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_322_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_323_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_323_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_324_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_324_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_325_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_325_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_326_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_326_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_327_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_327_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_328_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_328_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_329_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_329_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_330_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_330_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_331_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_331_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_332_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_332_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_333_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_333_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_334_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4097) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_334_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_335_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4099) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_335_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_336_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_336_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_337_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_337_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_338_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_338_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_339_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_339_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_340_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_340_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_341_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_341_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_342_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_342_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_343_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_343_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_344_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_344_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_345_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_345_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_346_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_346_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_347_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_347_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_348_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_348_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_349_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_349_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_350_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4117) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_350_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_351_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_4119) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_351_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_352_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_352_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_353_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_353_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_354_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_354_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_355_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_355_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_356_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_356_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_357_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_357_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_358_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_358_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_359_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_359_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_360_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_360_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_361_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_361_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_362_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_362_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_363_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_363_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_364_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_364_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_365_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_365_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_366_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_3964) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_366_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_367_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_3969) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_367_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_368_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_368_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_369_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4174 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_369_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_370_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_370_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_371_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4178 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_371_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_372_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_372_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_373_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4182 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_373_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_374_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_374_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_375_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4185 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_375_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_376_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_376_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_377_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4188 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_377_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_378_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_378_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_379_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4191 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_379_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_380_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_380_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_381_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4194 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_381_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_382_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_3988) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_382_reg <= z_out_5_19_4[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_383_reg <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[9])) | or_dcpl_4198 | or_dcpl_3990) ) begin
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_383_reg <= z_out_5_19_4[10:0];
    end
  end
  assign and_655_nl = (~((nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[1])
      ^ (nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[0]))) & (fsm_output[13]);
  assign and_661_nl = or_dcpl_2015 & (fsm_output[13]);
  assign and_667_nl = or_dcpl_2016 & (fsm_output[13]);
  assign Product2_1_jj_mux_nl = MUX_v_2_2_2((z_out[1:0]), (Accum1_ii_3_0_sva[1:0]),
      fsm_output[14]);
  assign nand_22_nl = ~(and_dcpl_2 & (~((fsm_output[9]) | (fsm_output[11]))));
  assign Product2_1_jj_Product2_1_jj_and_nl = MUX_v_2_2_2(2'b00, Product2_1_jj_mux_nl,
      nand_22_nl);
  assign Product1_ii_Product1_ii_mux_nl = MUX_v_4_2_2(z_out, ({2'b00 , Product2_1_jj_Product2_1_jj_and_nl}),
      Accum1_ii_3_0_sva_mx0c3);
  assign Accum1_ii_not_1_nl = ~ Accum1_ii_3_0_sva_mx0c0;
  assign Product1_mux_nl = MUX_v_16_14_2((input_1_rsci_idat[15:0]), (input_1_rsci_idat[31:16]),
      (input_1_rsci_idat[47:32]), (input_1_rsci_idat[63:48]), (input_1_rsci_idat[79:64]),
      (input_1_rsci_idat[95:80]), (input_1_rsci_idat[111:96]), (input_1_rsci_idat[127:112]),
      (input_1_rsci_idat[143:128]), (input_1_rsci_idat[159:144]), (input_1_rsci_idat[175:160]),
      (input_1_rsci_idat[191:176]), (input_1_rsci_idat[207:192]), (input_1_rsci_idat[223:208]),
      Accum1_ii_3_0_sva);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_or_nl = and_5052_rgt | and_5057_rgt;
  assign nor_23_nl = ~(((~((fsm_output[12]) | (fsm_output[7]))) & (~((fsm_output[4])
      | (fsm_output[10]))) & (~((fsm_output[11]) | (fsm_output[2]) | (fsm_output[6]))))
      | and_5035_cse);
  assign Product2_jj_and_nl = MUX_v_7_2_2(7'b0000000, (z_out_2[6:0]), nor_23_nl);
  assign or_7339_nl = (fsm_output[7]) | (fsm_output[6]) | (fsm_output[11]) | ((~
      Result_and_1_tmp) & (fsm_output[10]));
  assign mux_nl = MUX_v_7_2_2(Product2_jj_and_nl, (Result_ires_7_0_sva_1[6:0]), or_7339_nl);
  assign and_5067_nl = and_dcpl_35 & and_dcpl_32 & (fsm_output[4]);
  assign and_5074_nl = and_dcpl_35 & and_dcpl_38 & (fsm_output[4]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_or_4_nl = and_5081_rgt |
      and_5086_rgt;
  assign and_5095_nl = and_dcpl_49 & and_dcpl_32 & (fsm_output[4]);
  assign and_5102_nl = and_dcpl_52 & and_dcpl_21 & (fsm_output[4]);
  assign and_5109_nl = and_dcpl_49 & and_dcpl_38 & (fsm_output[4]);
  assign and_5116_nl = and_dcpl_52 & and_dcpl_41 & (fsm_output[4]);
  assign and_5123_nl = and_dcpl_35 & and_dcpl_56 & (fsm_output[4]);
  assign and_5130_nl = and_dcpl_24 & and_dcpl_58 & (fsm_output[4]);
  assign and_5137_nl = and_dcpl_35 & and_dcpl_60 & (fsm_output[4]);
  assign and_5144_nl = and_dcpl_24 & and_dcpl_62 & (fsm_output[4]);
  assign and_5151_nl = and_dcpl_49 & and_dcpl_56 & (fsm_output[4]);
  assign and_5158_nl = and_dcpl_52 & and_dcpl_58 & (fsm_output[4]);
  assign and_5165_nl = and_dcpl_49 & and_dcpl_60 & (fsm_output[4]);
  assign and_5172_nl = and_dcpl_52 & and_dcpl_62 & (fsm_output[4]);
  assign and_5179_nl = and_dcpl_35 & and_dcpl_62 & (fsm_output[4]);
  assign and_5186_nl = and_dcpl_24 & and_dcpl_60 & (fsm_output[4]);
  assign and_5193_nl = and_dcpl_35 & and_dcpl_58 & (fsm_output[4]);
  assign and_5200_nl = and_dcpl_24 & and_dcpl_56 & (fsm_output[4]);
  assign and_5207_nl = and_dcpl_49 & and_dcpl_62 & (fsm_output[4]);
  assign nnet_dense_latency_input_t_layer2_t_config2_acc_or_23_nl = and_5214_rgt
      | and_5219_rgt;
  assign and_5228_nl = and_dcpl_49 & and_dcpl_58 & (fsm_output[4]);
  assign and_5235_nl = and_dcpl_52 & and_dcpl_56 & (fsm_output[4]);
  assign and_5242_nl = and_dcpl_35 & and_dcpl_41 & (fsm_output[4]);
  assign and_5249_nl = and_dcpl_24 & and_dcpl_38 & (fsm_output[4]);
  assign and_5256_nl = and_dcpl_35 & and_dcpl_21 & (fsm_output[4]);
  assign and_5263_nl = and_dcpl_24 & and_dcpl_32 & (fsm_output[4]);
  assign and_5270_nl = and_dcpl_49 & and_dcpl_41 & (fsm_output[4]);
  assign and_5277_nl = and_dcpl_52 & and_dcpl_38 & (fsm_output[4]);
  assign and_5284_nl = and_dcpl_49 & and_dcpl_21 & (fsm_output[4]);
  assign and_5291_nl = and_dcpl_52 & and_dcpl_32 & (fsm_output[4]);
  assign and_5298_nl = and_dcpl_86 & and_dcpl_32 & (fsm_output[4]);
  assign and_5305_nl = and_dcpl_89 & and_dcpl_21 & (fsm_output[4]);
  assign and_5319_nl = and_dcpl_89 & and_dcpl_41 & (fsm_output[4]);
  assign and_5333_nl = and_dcpl_95 & and_dcpl_21 & (fsm_output[4]);
  assign and_5340_nl = and_dcpl_93 & and_dcpl_38 & (fsm_output[4]);
  assign and_5354_nl = and_dcpl_86 & and_dcpl_56 & (fsm_output[4]);
  assign and_5361_nl = and_dcpl_89 & and_dcpl_58 & (fsm_output[4]);
  assign and_5368_nl = and_dcpl_86 & and_dcpl_60 & (fsm_output[4]);
  assign and_5375_nl = and_dcpl_89 & and_dcpl_62 & (fsm_output[4]);
  assign and_5382_nl = and_dcpl_93 & and_dcpl_56 & (fsm_output[4]);
  assign and_5389_nl = and_dcpl_95 & and_dcpl_58 & (fsm_output[4]);
  assign and_5396_nl = and_dcpl_93 & and_dcpl_60 & (fsm_output[4]);
  assign and_5403_nl = and_dcpl_95 & and_dcpl_62 & (fsm_output[4]);
  assign and_5410_nl = and_dcpl_86 & and_dcpl_62 & (fsm_output[4]);
  assign and_5417_nl = and_dcpl_89 & and_dcpl_60 & (fsm_output[4]);
  assign and_5424_nl = and_dcpl_86 & and_dcpl_58 & (fsm_output[4]);
  assign and_5431_nl = and_dcpl_89 & and_dcpl_56 & (fsm_output[4]);
  assign and_5438_nl = and_dcpl_93 & and_dcpl_62 & (fsm_output[4]);
  assign and_5445_nl = and_dcpl_95 & and_dcpl_60 & (fsm_output[4]);
  assign and_5452_nl = and_dcpl_93 & and_dcpl_58 & (fsm_output[4]);
  assign and_5461_nl = and_dcpl_95 & and_dcpl_56 & (fsm_output[4]);
  assign and_5468_nl = and_dcpl_86 & and_dcpl_41 & (fsm_output[4]);
  assign and_5475_nl = and_dcpl_89 & and_dcpl_38 & (fsm_output[4]);
  assign and_5482_nl = and_dcpl_86 & and_dcpl_21 & (fsm_output[4]);
  assign and_5489_nl = and_dcpl_89 & and_dcpl_32 & (fsm_output[4]);
  assign and_5496_nl = and_dcpl_93 & and_dcpl_41 & (fsm_output[4]);
  assign and_5503_nl = and_dcpl_95 & and_dcpl_38 & (fsm_output[4]);
  assign and_5510_nl = and_dcpl_93 & and_dcpl_21 & (fsm_output[4]);
  assign and_5517_nl = and_dcpl_95 & and_dcpl_32 & (fsm_output[4]);
  assign and_5524_nl = and_dcpl_123 & and_dcpl_32 & (fsm_output[4]);
  assign and_5531_nl = and_dcpl_125 & and_dcpl_21 & (fsm_output[4]);
  assign and_5538_nl = and_dcpl_123 & and_dcpl_38 & (fsm_output[4]);
  assign and_5545_nl = and_dcpl_125 & and_dcpl_41 & (fsm_output[4]);
  assign and_5552_nl = and_dcpl_129 & and_dcpl_32 & (fsm_output[4]);
  assign and_5559_nl = and_dcpl_131 & and_dcpl_21 & (fsm_output[4]);
  assign and_5566_nl = and_dcpl_129 & and_dcpl_38 & (fsm_output[4]);
  assign and_5580_nl = and_dcpl_123 & and_dcpl_56 & (fsm_output[4]);
  assign and_5587_nl = and_dcpl_125 & and_dcpl_58 & (fsm_output[4]);
  assign and_5594_nl = and_dcpl_123 & and_dcpl_60 & (fsm_output[4]);
  assign and_5601_nl = and_dcpl_125 & and_dcpl_62 & (fsm_output[4]);
  assign and_5608_nl = and_dcpl_129 & and_dcpl_56 & (fsm_output[4]);
  assign and_5615_nl = and_dcpl_131 & and_dcpl_58 & (fsm_output[4]);
  assign and_5629_nl = and_dcpl_131 & and_dcpl_62 & (fsm_output[4]);
  assign and_5636_nl = and_dcpl_123 & and_dcpl_62 & (fsm_output[4]);
  assign and_5643_nl = and_dcpl_125 & and_dcpl_60 & (fsm_output[4]);
  assign and_5650_nl = and_dcpl_123 & and_dcpl_58 & (fsm_output[4]);
  assign and_5657_nl = and_dcpl_125 & and_dcpl_56 & (fsm_output[4]);
  assign and_5664_nl = and_dcpl_129 & and_dcpl_62 & (fsm_output[4]);
  assign and_5671_nl = and_dcpl_131 & and_dcpl_60 & (fsm_output[4]);
  assign and_5678_nl = and_dcpl_129 & and_dcpl_58 & (fsm_output[4]);
  assign and_5685_nl = and_dcpl_131 & and_dcpl_56 & (fsm_output[4]);
  assign and_5692_nl = and_dcpl_123 & and_dcpl_41 & (fsm_output[4]);
  assign and_5699_nl = and_dcpl_125 & and_dcpl_38 & (fsm_output[4]);
  assign and_5706_nl = and_dcpl_123 & and_dcpl_21 & (fsm_output[4]);
  assign and_5713_nl = and_dcpl_125 & and_dcpl_32 & (fsm_output[4]);
  assign and_5720_nl = and_dcpl_129 & and_dcpl_41 & (fsm_output[4]);
  assign and_5727_nl = and_dcpl_131 & and_dcpl_38 & (fsm_output[4]);
  assign and_5734_nl = and_dcpl_129 & and_dcpl_21 & (fsm_output[4]);
  assign and_5741_nl = and_dcpl_131 & and_dcpl_32 & (fsm_output[4]);
  assign and_5748_nl = and_dcpl_159 & and_dcpl_32 & (fsm_output[4]);
  assign and_5755_nl = and_dcpl_161 & and_dcpl_21 & (fsm_output[4]);
  assign and_5769_nl = and_dcpl_161 & and_dcpl_41 & (fsm_output[4]);
  assign and_5776_nl = and_dcpl_165 & and_dcpl_32 & (fsm_output[4]);
  assign and_5783_nl = and_dcpl_167 & and_dcpl_21 & (fsm_output[4]);
  assign and_5790_nl = and_dcpl_165 & and_dcpl_38 & (fsm_output[4]);
  assign and_5797_nl = and_dcpl_167 & and_dcpl_41 & (fsm_output[4]);
  assign and_5804_nl = and_dcpl_159 & and_dcpl_56 & (fsm_output[4]);
  assign and_5811_nl = and_dcpl_161 & and_dcpl_58 & (fsm_output[4]);
  assign and_5818_nl = and_dcpl_159 & and_dcpl_60 & (fsm_output[4]);
  assign and_5825_nl = and_dcpl_161 & and_dcpl_62 & (fsm_output[4]);
  assign and_5832_nl = and_dcpl_165 & and_dcpl_56 & (fsm_output[4]);
  assign and_5839_nl = and_dcpl_167 & and_dcpl_58 & (fsm_output[4]);
  assign and_5846_nl = and_dcpl_165 & and_dcpl_60 & (fsm_output[4]);
  assign and_5853_nl = and_dcpl_167 & and_dcpl_62 & (fsm_output[4]);
  assign and_5860_nl = and_dcpl_159 & and_dcpl_62 & (fsm_output[4]);
  assign and_5867_nl = and_dcpl_161 & and_dcpl_60 & (fsm_output[4]);
  assign and_5874_nl = and_dcpl_159 & and_dcpl_58 & (fsm_output[4]);
  assign and_5881_nl = and_dcpl_161 & and_dcpl_56 & (fsm_output[4]);
  assign and_5888_nl = and_dcpl_165 & and_dcpl_62 & (fsm_output[4]);
  assign and_5895_nl = and_dcpl_167 & and_dcpl_60 & (fsm_output[4]);
  assign and_5902_nl = and_dcpl_165 & and_dcpl_58 & (fsm_output[4]);
  assign and_5909_nl = and_dcpl_167 & and_dcpl_56 & (fsm_output[4]);
  assign and_5916_nl = and_dcpl_159 & and_dcpl_41 & (fsm_output[4]);
  assign and_5923_nl = and_dcpl_161 & and_dcpl_38 & (fsm_output[4]);
  assign and_5930_nl = and_dcpl_159 & and_dcpl_21 & (fsm_output[4]);
  assign and_5937_nl = and_dcpl_161 & and_dcpl_32 & (fsm_output[4]);
  assign and_5944_nl = and_dcpl_165 & and_dcpl_41 & (fsm_output[4]);
  assign and_5951_nl = and_dcpl_167 & and_dcpl_38 & (fsm_output[4]);
  assign and_5958_nl = and_dcpl_165 & and_dcpl_21 & (fsm_output[4]);
  assign or_7335_nl = (fsm_output[10]) | (fsm_output[6]);
  assign and_nl = MUX_v_7_2_2(7'b0000000, (nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[6:0]),
      or_7335_nl);
  assign Product2_1_jj_mux_1_nl = MUX_v_2_2_2((z_out_1[1:0]), (nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[1:0]),
      fsm_output[14]);
  assign not_568_nl = ~ and_dcpl_2;
  assign Product2_1_jj_Product2_1_jj_and_1_nl = MUX_v_2_2_2(2'b00, Product2_1_jj_mux_1_nl,
      not_568_nl);
  assign Product2_jj_Product2_jj_and_1_nl = MUX_v_7_2_2(7'b0000000, (nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_7_0_sva_1[6:0]),
      (fsm_output[10]));
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((Accum2_mux_131[8:1]), 8'b11111111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1);
  assign Product1_mux_3_nl = MUX_v_2_2_2((Accum1_ii_3_0_sva[3:2]), (signext_2_1(Accum1_ii_3_0_sva[1])),
      or_7342_cse);
  assign nl_z_out = ({Product1_mux_3_nl , (Accum1_ii_3_0_sva[1:0])}) + 4'b0001;
  assign z_out = nl_z_out[3:0];
  assign or_7367_nl = (fsm_output[5]) | (fsm_output[3]);
  assign nnet_linear_layer5_t_result_t_linear_config6_for_mux_5_nl = MUX_v_4_2_2((signext_4_2(nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[1:0])),
      ({1'b1 , (z_out[3:1])}), or_7367_nl);
  assign nl_z_out_1 = nnet_linear_layer5_t_result_t_linear_config6_for_mux_5_nl +
      4'b0001;
  assign z_out_1 = nl_z_out_1[3:0];
  assign or_7368_nl = (fsm_output[12]) | (fsm_output[8]) | (fsm_output[4]) | (fsm_output[2]);
  assign nnet_linear_layer2_t_layer3_t_linear_config3_for_mux1h_1_nl = MUX1HOT_v_7_5_2((nnet_linear_layer2_t_layer3_t_linear_config3_for_ii_7_0_sva_1[6:0]),
      (nnet_relu_layer3_t_layer4_t_relu_config4_for_ii_7_0_sva_1[6:0]), (Result_ires_7_0_sva_1[6:0]),
      Product1_1_ii_7_0_sva_6_0, ({5'b11111 , (z_out[1:0])}), {(fsm_output[7]) ,
      (fsm_output[6]) , or_7368_nl , (fsm_output[10]) , or_7342_cse});
  assign nl_z_out_2 = conv_u2u_7_8(nnet_linear_layer2_t_layer3_t_linear_config3_for_mux1h_1_nl)
      + 8'b00000001;
  assign z_out_2 = nl_z_out_2[7:0];
  assign nl_Product2_1_index_acc_sdt = conv_u2u_7_8(Product2_1_index_mux_cse) + conv_u2u_2_8(Accum1_ii_3_0_sva[1:0]);
  assign Product2_1_index_acc_sdt = nl_Product2_1_index_acc_sdt[7:0];
  assign nl_z_out_4_8_1 = conv_u2u_7_8(Product2_1_index_acc_sdt[7:1]) + conv_u2u_7_8(Product2_1_index_mux_cse);
  assign z_out_4_8_1 = nl_z_out_4_8_1[7:0];
  assign nnet_product_mult_input_t_config2_weight_t_product_mux_2_nl = MUX_v_5_2_2(ROM_1i11_1o5_815f6a3dbd0daa2d77beb65dd6cecbbc31_1,
      ROM_1i9_1o5_4a143e9cb1f27bd26e0331874cec74ad2f_1, fsm_output[9]);
  assign nnet_product_mult_input_t_config2_weight_t_product_mux_3_nl = MUX_v_16_2_2(nnet_dense_latency_input_t_layer2_t_config2_acc_0_lpi_3,
      ({6'b000000 , layer4_out_9_lpi_2_dfm , layer4_out_8_1_lpi_2_dfm , layer4_out_0_lpi_2_dfm}),
      fsm_output[9]);
  assign nl_mul_nl = $signed(nnet_product_mult_input_t_config2_weight_t_product_mux_2_nl)
      * $signed(nnet_product_mult_input_t_config2_weight_t_product_mux_3_nl);
  assign mul_nl = nl_mul_nl[19:0];
  assign z_out_5_19_4 = readslicef_20_16_4(mul_nl);
  assign Accum2_mux_133_nl = MUX_v_16_2_2(Accum2_mux_131, Accum2_1_mux_6, fsm_output[11]);
  assign Accum2_mux_135_nl = MUX_v_16_1792_2(nnet_dense_latency_input_t_layer2_t_config2_mult_0_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_2_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_3_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_4_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_5_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_6_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_7_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_8_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_9_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_10_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_11_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_12_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_13_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_14_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_15_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_16_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_17_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_18_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_19_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_20_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_21_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_22_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_23_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_24_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_25_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_26_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_27_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_28_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_29_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_30_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_31_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_32_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_33_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_34_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_35_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_36_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_37_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_38_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_39_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_40_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_41_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_42_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_43_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_44_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_45_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_46_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_47_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_48_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_49_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_50_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_51_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_52_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_53_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_54_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_55_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_56_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_57_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_58_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_59_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_60_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_61_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_62_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_63_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_64_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_65_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_66_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_67_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_68_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_69_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_70_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_71_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_72_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_73_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_74_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_75_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_76_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_77_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_78_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_79_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_80_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_81_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_82_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_83_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_84_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_85_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_86_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_87_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_88_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_89_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_90_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_91_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_92_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_93_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_94_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_95_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_96_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_97_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_98_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_99_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_100_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_101_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_102_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_103_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_104_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_105_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_106_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_107_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_108_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_109_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_110_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_111_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_112_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_113_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_114_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_115_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_116_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_117_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_118_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_119_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_120_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_121_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_122_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_123_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_124_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_125_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_126_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_127_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_128_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_129_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_130_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_131_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_132_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_133_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_134_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_135_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_136_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_137_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_138_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_139_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_140_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_141_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_142_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_143_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_144_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_145_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_146_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_147_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_148_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_149_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_150_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_151_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_152_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_153_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_154_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_155_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_156_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_157_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_158_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_159_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_160_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_161_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_162_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_163_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_164_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_165_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_166_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_167_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_168_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_169_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_170_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_171_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_172_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_173_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_174_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_175_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_176_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_177_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_178_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_179_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_180_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_181_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_182_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_183_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_184_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_185_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_186_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_187_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_188_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_189_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_190_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_191_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_192_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_193_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_194_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_195_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_196_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_197_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_198_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_199_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_200_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_201_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_202_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_203_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_204_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_205_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_206_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_207_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_208_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_209_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_210_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_211_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_212_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_213_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_214_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_215_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_216_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_217_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_218_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_219_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_220_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_221_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_222_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_223_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_224_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_225_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_226_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_227_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_228_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_229_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_230_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_231_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_232_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_233_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_234_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_235_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_236_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_237_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_238_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_239_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_240_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_241_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_242_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_243_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_244_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_245_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_246_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_247_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_248_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_249_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_250_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_251_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_252_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_253_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_254_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_255_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_256_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_257_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_258_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_259_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_260_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_261_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_262_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_263_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_264_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_265_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_266_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_267_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_268_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_269_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_270_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_271_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_272_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_273_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_274_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_275_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_276_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_277_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_278_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_279_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_280_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_281_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_282_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_283_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_284_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_285_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_286_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_287_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_288_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_289_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_290_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_291_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_292_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_293_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_294_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_295_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_296_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_297_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_298_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_299_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_300_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_301_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_302_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_303_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_304_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_305_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_306_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_307_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_308_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_309_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_310_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_311_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_312_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_313_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_314_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_315_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_316_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_317_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_318_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_319_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_320_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_321_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_322_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_323_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_324_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_325_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_326_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_327_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_328_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_329_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_330_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_331_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_332_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_333_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_334_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_335_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_336_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_337_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_338_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_339_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_340_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_341_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_342_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_343_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_344_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_345_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_346_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_347_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_348_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_349_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_350_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_351_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_352_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_353_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_354_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_355_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_356_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_357_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_358_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_359_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_360_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_361_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_362_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_363_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_364_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_365_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_366_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_367_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_368_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_369_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_370_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_371_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_372_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_373_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_374_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_375_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_376_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_377_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_378_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_379_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_380_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_381_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_382_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_383_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_384_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_385_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_386_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_387_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_388_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_389_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_390_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_391_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_392_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_393_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_394_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_395_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_396_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_397_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_398_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_399_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_400_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_401_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_402_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_403_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_404_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_405_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_406_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_407_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_408_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_409_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_410_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_411_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_412_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_413_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_414_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_415_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_416_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_417_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_418_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_419_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_420_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_421_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_422_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_423_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_424_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_425_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_426_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_427_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_428_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_429_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_430_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_431_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_432_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_433_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_434_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_435_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_436_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_437_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_438_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_439_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_440_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_441_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_442_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_443_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_444_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_445_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_446_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_447_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_448_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_449_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_450_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_451_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_452_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_453_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_454_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_455_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_456_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_457_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_458_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_459_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_460_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_461_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_462_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_463_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_464_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_465_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_466_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_467_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_468_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_469_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_470_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_471_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_472_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_473_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_474_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_475_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_476_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_477_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_478_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_479_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_480_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_481_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_482_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_483_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_484_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_485_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_486_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_487_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_488_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_489_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_490_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_491_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_492_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_493_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_494_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_495_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_496_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_497_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_498_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_499_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_500_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_501_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_502_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_503_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_504_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_505_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_506_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_507_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_508_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_509_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_510_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_511_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_512_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_513_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_514_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_515_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_516_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_517_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_518_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_519_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_520_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_521_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_522_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_523_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_524_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_525_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_526_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_527_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_528_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_529_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_530_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_531_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_532_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_533_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_534_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_535_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_536_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_537_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_538_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_539_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_540_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_541_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_542_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_543_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_544_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_545_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_546_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_547_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_548_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_549_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_550_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_551_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_552_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_553_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_554_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_555_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_556_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_557_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_558_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_559_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_560_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_561_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_562_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_563_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_564_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_565_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_566_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_567_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_568_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_569_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_570_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_571_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_572_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_573_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_574_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_575_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_576_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_577_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_578_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_579_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_580_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_581_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_582_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_583_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_584_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_585_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_586_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_587_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_588_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_589_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_590_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_591_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_592_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_593_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_594_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_595_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_596_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_597_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_598_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_599_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_600_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_601_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_602_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_603_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_604_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_605_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_606_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_607_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_608_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_609_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_610_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_611_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_612_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_613_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_614_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_615_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_616_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_617_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_618_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_619_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_620_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_621_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_622_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_623_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_624_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_625_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_626_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_627_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_628_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_629_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_630_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_631_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_632_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_633_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_634_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_635_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_636_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_637_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_638_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_639_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_640_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_641_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_642_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_643_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_644_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_645_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_646_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_647_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_648_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_649_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_650_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_651_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_652_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_653_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_654_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_655_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_656_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_657_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_658_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_659_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_660_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_661_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_662_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_663_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_664_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_665_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_666_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_667_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_668_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_669_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_670_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_671_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_672_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_673_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_674_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_675_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_676_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_677_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_678_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_679_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_680_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_681_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_682_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_683_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_684_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_685_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_686_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_687_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_688_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_689_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_690_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_691_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_692_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_693_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_694_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_695_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_696_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_697_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_698_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_699_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_700_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_701_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_702_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_703_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_704_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_705_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_706_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_707_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_708_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_709_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_710_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_711_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_712_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_713_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_714_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_715_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_716_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_717_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_718_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_719_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_720_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_721_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_722_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_723_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_724_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_725_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_726_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_727_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_728_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_729_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_730_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_731_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_732_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_733_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_734_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_735_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_736_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_737_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_738_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_739_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_740_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_741_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_742_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_743_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_744_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_745_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_746_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_747_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_748_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_749_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_750_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_751_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_752_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_753_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_754_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_755_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_756_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_757_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_758_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_759_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_760_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_761_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_762_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_763_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_764_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_765_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_766_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_767_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_768_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_769_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_770_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_771_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_772_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_773_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_774_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_775_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_776_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_777_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_778_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_779_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_780_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_781_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_782_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_783_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_784_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_785_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_786_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_787_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_788_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_789_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_790_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_791_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_792_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_793_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_794_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_795_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_796_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_797_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_798_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_799_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_800_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_801_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_802_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_803_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_804_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_805_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_806_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_807_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_808_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_809_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_810_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_811_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_812_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_813_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_814_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_815_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_816_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_817_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_818_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_819_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_820_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_821_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_822_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_823_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_824_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_825_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_826_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_827_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_828_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_829_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_830_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_831_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_832_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_833_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_834_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_835_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_836_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_837_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_838_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_839_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_840_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_841_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_842_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_843_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_844_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_845_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_846_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_847_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_848_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_849_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_850_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_851_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_852_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_853_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_854_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_855_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_856_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_857_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_858_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_859_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_860_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_861_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_862_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_863_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_864_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_865_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_866_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_867_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_868_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_869_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_870_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_871_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_872_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_873_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_874_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_875_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_876_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_877_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_878_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_879_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_880_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_881_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_882_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_883_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_884_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_885_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_886_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_887_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_888_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_889_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_890_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_891_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_892_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_893_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_894_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_895_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_896_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_897_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_898_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_899_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_900_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_901_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_902_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_903_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_904_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_905_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_906_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_907_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_908_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_909_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_910_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_911_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_912_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_913_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_914_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_915_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_916_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_917_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_918_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_919_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_920_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_921_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_922_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_923_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_924_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_925_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_926_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_927_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_928_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_929_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_930_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_931_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_932_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_933_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_934_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_935_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_936_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_937_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_938_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_939_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_940_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_941_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_942_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_943_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_944_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_945_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_946_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_947_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_948_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_949_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_950_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_951_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_952_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_953_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_954_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_955_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_956_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_957_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_958_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_959_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_960_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_961_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_962_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_963_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_964_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_965_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_966_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_967_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_968_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_969_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_970_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_971_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_972_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_973_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_974_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_975_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_976_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_977_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_978_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_979_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_980_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_981_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_982_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_983_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_984_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_985_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_986_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_987_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_988_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_989_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_990_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_991_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_992_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_993_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_994_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_995_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_996_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_997_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_998_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_999_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1000_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1001_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1002_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1003_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1004_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1005_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1006_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1007_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1008_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1009_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1010_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1011_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1012_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1013_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1014_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1015_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1016_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1017_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1018_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1019_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1020_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1021_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1022_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1023_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1024_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1025_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1026_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1027_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1028_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1029_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1030_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1031_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1032_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1033_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1034_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1035_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1036_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1037_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1038_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1039_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1040_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1041_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1042_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1043_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1044_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1045_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1046_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1047_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1048_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1049_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1050_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1051_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1052_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1053_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1054_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1055_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1056_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1057_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1058_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1059_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1060_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1061_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1062_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1063_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1064_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1065_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1066_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1067_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1068_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1069_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1070_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1071_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1072_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1073_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1074_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1075_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1076_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1077_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1078_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1079_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1080_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1081_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1082_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1083_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1084_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1085_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1086_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1087_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1088_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1089_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1090_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1091_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1092_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1093_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1094_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1095_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1096_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1097_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1098_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1099_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1100_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1101_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1102_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1103_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1104_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1105_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1106_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1107_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1108_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1109_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1110_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1111_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1112_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1113_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1114_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1115_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1116_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1117_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1118_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1119_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1120_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1121_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1122_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1123_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1124_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1125_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1126_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1127_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1128_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1129_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1130_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1131_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1132_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1133_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1134_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1135_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1136_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1137_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1138_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1139_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1140_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1141_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1142_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1143_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1144_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1145_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1146_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1147_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1148_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1149_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1150_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1151_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1152_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1153_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1154_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1155_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1156_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1157_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1158_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1159_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1160_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1161_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1162_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1163_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1164_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1165_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1166_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1167_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1168_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1169_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1170_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1171_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1172_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1173_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1174_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1175_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1176_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1177_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1178_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1179_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1180_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1181_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1182_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1183_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1184_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1185_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1186_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1187_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1188_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1189_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1190_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1191_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1192_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1193_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1194_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1195_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1196_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1197_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1198_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1199_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1200_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1201_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1202_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1203_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1204_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1205_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1206_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1207_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1208_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1209_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1210_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1211_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1212_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1213_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1214_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1215_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1216_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1217_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1218_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1219_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1220_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1221_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1222_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1223_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1224_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1225_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1226_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1227_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1228_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1229_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1230_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1231_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1232_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1233_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1234_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1235_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1236_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1237_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1238_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1239_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1240_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1241_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1242_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1243_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1244_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1245_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1246_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1247_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1248_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1249_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1250_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1251_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1252_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1253_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1254_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1255_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1256_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1257_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1258_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1259_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1260_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1261_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1262_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1263_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1264_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1265_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1266_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1267_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1268_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1269_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1270_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1271_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1272_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1273_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1274_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1275_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1276_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1277_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1278_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1279_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1280_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1281_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1282_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1283_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1284_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1285_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1286_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1287_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1288_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1289_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1290_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1291_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1292_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1293_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1294_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1295_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1296_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1297_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1298_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1299_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1300_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1301_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1302_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1303_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1304_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1305_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1306_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1307_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1308_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1309_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1310_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1311_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1312_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1313_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1314_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1315_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1316_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1317_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1318_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1319_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1320_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1321_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1322_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1323_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1324_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1325_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1326_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1327_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1328_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1329_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1330_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1331_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1332_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1333_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1334_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1335_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1336_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1337_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1338_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1339_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1340_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1341_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1342_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1343_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1344_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1345_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1346_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1347_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1348_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1349_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1350_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1351_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1352_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1353_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1354_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1355_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1356_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1357_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1358_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1359_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1360_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1361_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1362_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1363_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1364_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1365_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1366_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1367_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1368_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1369_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1370_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1371_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1372_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1373_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1374_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1375_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1376_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1377_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1378_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1379_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1380_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1381_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1382_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1383_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1384_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1385_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1386_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1387_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1388_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1389_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1390_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1391_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1392_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1393_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1394_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1395_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1396_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1397_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1398_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1399_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1400_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1401_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1402_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1403_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1404_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1405_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1406_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1407_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1408_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1409_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1410_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1411_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1412_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1413_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1414_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1415_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1416_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1417_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1418_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1419_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1420_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1421_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1422_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1423_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1424_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1425_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1426_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1427_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1428_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1429_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1430_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1431_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1432_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1433_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1434_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1435_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1436_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1437_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1438_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1439_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1440_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1441_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1442_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1443_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1444_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1445_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1446_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1447_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1448_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1449_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1450_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1451_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1452_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1453_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1454_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1455_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1456_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1457_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1458_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1459_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1460_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1461_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1462_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1463_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1464_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1465_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1466_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1467_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1468_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1469_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1470_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1471_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1472_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1473_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1474_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1475_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1476_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1477_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1478_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1479_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1480_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1481_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1482_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1483_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1484_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1485_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1486_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1487_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1488_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1489_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1490_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1491_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1492_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1493_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1494_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1495_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1496_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1497_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1498_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1499_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1500_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1501_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1502_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1503_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1504_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1505_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1506_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1507_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1508_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1509_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1510_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1511_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1512_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1513_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1514_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1515_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1516_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1517_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1518_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1519_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1520_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1521_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1522_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1523_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1524_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1525_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1526_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1527_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1528_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1529_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1530_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1531_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1532_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1533_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1534_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1535_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1536_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1537_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1538_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1539_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1540_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1541_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1542_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1543_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1544_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1545_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1546_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1547_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1548_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1549_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1550_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1551_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1552_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1553_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1554_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1555_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1556_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1557_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1558_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1559_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1560_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1561_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1562_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1563_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1564_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1565_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1566_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1567_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1568_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1569_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1570_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1571_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1572_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1573_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1574_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1575_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1576_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1577_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1578_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1579_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1580_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1581_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1582_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1583_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1584_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1585_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1586_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1587_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1588_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1589_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1590_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1591_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1592_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1593_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1594_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1595_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1596_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1597_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1598_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1599_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1600_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1601_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1602_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1603_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1604_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1605_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1606_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1607_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1608_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1609_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1610_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1611_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1612_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1613_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1614_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1615_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1616_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1617_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1618_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1619_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1620_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1621_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1622_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1623_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1624_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1625_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1626_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1627_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1628_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1629_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1630_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1631_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1632_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1633_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1634_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1635_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1636_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1637_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1638_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1639_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1640_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1641_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1642_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1643_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1644_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1645_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1646_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1647_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1648_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1649_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1650_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1651_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1652_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1653_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1654_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1655_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1656_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1657_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1658_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1659_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1660_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1661_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1662_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1663_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1664_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1665_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1666_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1667_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1668_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1669_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1670_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1671_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1672_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1673_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1674_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1675_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1676_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1677_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1678_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1679_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1680_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1681_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1682_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1683_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1684_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1685_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1686_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1687_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1688_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1689_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1690_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1691_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1692_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1693_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1694_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1695_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1696_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1697_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1698_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1699_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1700_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1701_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1702_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1703_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1704_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1705_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1706_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1707_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1708_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1709_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1710_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1711_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1712_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1713_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1714_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1715_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1716_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1717_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1718_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1719_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1720_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1721_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1722_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1723_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1724_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1725_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1726_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1727_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1728_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1729_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1730_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1731_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1732_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1733_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1734_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1735_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1736_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1737_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1738_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1739_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1740_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1741_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1742_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1743_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1744_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1745_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1746_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1747_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1748_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1749_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1750_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1751_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1752_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1753_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1754_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1755_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1756_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1757_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1758_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1759_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1760_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1761_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1762_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1763_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1764_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1765_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1766_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1767_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1768_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1769_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1770_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1771_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1772_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1773_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1774_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1775_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1776_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1777_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1778_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1779_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1780_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1781_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1782_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1783_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1784_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1785_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1786_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1787_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1788_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1789_lpi_3, nnet_dense_latency_input_t_layer2_t_config2_mult_1790_lpi_3,
      nnet_dense_latency_input_t_layer2_t_config2_mult_1791_lpi_3, {Accum1_ii_3_0_sva
      , (Result_ires_7_0_sva_1[6:0])});
  assign Accum2_1_mux_7_nl = MUX_v_16_384_2(({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_0_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_0_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_1_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_1_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_2_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_2_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_3_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_3_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_4_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_4_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_5_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_5_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_6_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_6_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_7_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_7_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_8_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_8_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_9_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_9_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_10_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_10_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_11_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_11_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_12_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_12_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_13_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_13_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_14_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_14_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_15_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_15_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_16_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_16_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_17_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_17_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_18_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_18_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_19_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_19_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_20_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_20_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_21_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_21_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_22_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_22_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_23_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_23_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_24_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_24_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_25_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_25_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_26_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_26_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_27_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_27_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_28_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_28_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_29_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_29_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_30_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_30_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_31_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_31_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_32_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_32_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_33_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_33_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_34_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_34_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_35_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_35_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_36_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_36_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_37_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_37_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_38_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_38_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_39_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_39_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_40_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_40_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_41_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_41_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_42_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_42_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_43_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_43_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_44_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_44_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_45_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_45_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_46_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_46_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_47_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_47_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_48_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_48_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_49_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_49_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_50_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_50_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_51_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_51_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_52_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_52_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_53_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_53_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_54_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_54_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_55_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_55_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_56_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_56_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_57_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_57_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_58_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_58_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_59_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_59_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_60_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_60_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_61_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_61_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_62_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_62_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_63_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_63_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_64_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_64_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_65_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_65_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_66_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_66_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_67_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_67_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_68_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_68_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_69_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_69_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_70_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_70_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_71_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_71_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_72_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_72_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_73_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_73_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_74_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_74_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_75_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_75_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_76_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_76_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_77_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_77_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_78_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_78_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_79_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_79_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_80_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_80_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_81_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_81_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_82_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_82_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_83_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_83_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_84_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_84_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_85_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_85_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_86_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_86_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_87_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_87_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_88_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_88_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_89_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_89_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_90_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_90_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_91_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_91_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_92_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_92_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_93_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_93_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_94_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_94_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_95_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_95_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_96_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_96_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_97_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_97_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_98_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_98_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_99_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_99_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_100_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_100_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_101_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_101_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_102_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_102_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_103_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_103_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_104_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_104_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_105_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_105_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_106_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_106_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_107_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_107_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_108_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_108_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_109_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_109_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_110_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_110_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_111_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_111_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_112_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_112_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_113_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_113_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_114_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_114_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_115_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_115_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_116_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_116_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_117_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_117_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_118_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_118_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_119_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_119_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_120_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_120_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_121_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_121_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_122_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_122_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_123_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_123_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_124_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_124_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_125_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_125_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_126_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_126_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_127_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_127_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_128_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_128_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_129_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_129_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_130_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_130_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_131_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_131_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_132_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_132_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_133_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_133_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_134_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_134_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_135_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_135_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_136_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_136_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_137_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_137_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_138_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_138_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_139_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_139_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_140_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_140_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_141_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_141_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_142_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_142_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_143_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_143_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_144_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_144_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_145_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_145_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_146_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_146_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_147_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_147_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_148_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_148_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_149_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_149_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_150_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_150_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_151_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_151_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_152_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_152_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_153_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_153_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_154_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_154_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_155_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_155_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_156_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_156_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_157_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_157_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_158_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_158_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_159_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_159_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_160_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_160_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_161_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_161_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_162_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_162_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_163_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_163_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_164_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_164_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_165_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_165_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_166_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_166_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_167_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_167_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_168_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_168_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_169_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_169_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_170_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_170_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_171_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_171_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_172_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_172_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_173_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_173_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_174_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_174_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_175_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_175_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_176_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_176_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_177_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_177_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_178_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_178_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_179_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_179_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_180_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_180_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_181_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_181_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_182_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_182_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_183_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_183_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_184_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_184_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_185_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_185_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_186_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_186_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_187_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_187_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_188_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_188_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_189_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_189_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_190_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_190_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_191_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_191_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_192_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_192_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_193_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_193_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_194_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_194_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_195_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_195_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_196_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_196_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_197_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_197_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_198_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_198_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_199_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_199_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_200_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_200_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_201_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_201_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_202_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_202_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_203_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_203_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_204_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_204_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_205_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_205_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_206_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_206_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_207_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_207_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_208_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_208_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_209_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_209_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_210_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_210_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_211_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_211_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_212_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_212_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_213_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_213_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_214_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_214_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_215_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_215_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_216_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_216_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_217_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_217_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_218_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_218_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_219_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_219_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_220_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_220_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_221_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_221_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_222_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_222_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_223_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_223_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_224_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_224_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_225_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_225_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_226_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_226_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_227_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_227_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_228_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_228_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_229_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_229_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_230_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_230_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_231_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_231_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_232_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_232_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_233_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_233_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_234_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_234_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_235_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_235_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_236_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_236_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_237_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_237_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_238_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_238_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_239_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_239_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_240_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_240_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_241_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_241_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_242_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_242_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_243_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_243_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_244_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_244_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_245_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_245_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_246_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_246_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_247_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_247_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_248_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_248_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_249_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_249_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_250_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_250_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_251_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_251_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_252_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_252_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_253_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_253_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_254_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_254_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_255_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_255_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_256_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_256_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_257_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_257_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_258_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_258_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_259_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_259_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_260_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_260_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_261_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_261_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_262_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_262_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_263_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_263_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_264_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_264_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_265_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_265_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_266_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_266_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_267_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_267_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_268_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_268_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_269_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_269_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_270_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_270_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_271_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_271_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_272_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_272_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_273_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_273_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_274_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_274_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_275_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_275_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_276_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_276_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_277_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_277_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_278_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_278_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_279_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_279_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_280_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_280_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_281_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_281_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_282_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_282_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_283_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_283_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_284_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_284_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_285_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_285_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_286_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_286_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_287_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_287_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_288_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_288_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_289_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_289_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_290_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_290_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_291_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_291_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_292_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_292_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_293_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_293_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_294_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_294_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_295_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_295_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_296_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_296_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_297_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_297_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_298_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_298_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_299_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_299_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_300_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_300_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_301_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_301_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_302_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_302_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_303_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_303_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_304_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_304_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_305_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_305_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_306_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_306_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_307_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_307_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_308_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_308_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_309_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_309_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_310_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_310_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_311_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_311_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_312_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_312_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_313_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_313_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_314_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_314_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_315_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_315_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_316_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_316_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_317_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_317_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_318_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_318_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_319_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_319_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_320_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_320_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_321_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_321_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_322_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_322_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_323_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_323_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_324_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_324_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_325_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_325_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_326_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_326_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_327_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_327_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_328_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_328_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_329_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_329_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_330_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_330_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_331_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_331_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_332_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_332_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_333_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_333_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_334_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_334_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_335_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_335_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_336_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_336_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_337_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_337_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_338_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_338_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_339_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_339_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_340_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_340_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_341_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_341_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_342_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_342_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_343_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_343_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_344_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_344_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_345_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_345_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_346_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_346_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_347_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_347_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_348_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_348_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_349_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_349_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_350_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_350_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_351_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_351_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_352_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_352_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_353_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_353_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_354_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_354_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_355_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_355_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_356_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_356_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_357_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_357_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_358_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_358_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_359_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_359_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_360_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_360_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_361_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_361_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_362_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_362_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_363_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_363_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_364_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_364_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_365_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_365_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_366_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_366_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_367_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_367_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_368_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_368_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_369_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_369_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_370_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_370_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_371_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_371_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_372_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_372_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_373_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_373_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_374_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_374_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_375_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_375_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_376_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_376_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_377_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_377_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_378_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_378_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_379_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_379_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_380_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_380_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_381_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_381_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_382_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_382_reg}), ({{5{reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_383_reg[10]}},
      reg_nnet_dense_latency_layer4_t_layer5_t_config5_mult_383_reg}), {z_out_4_8_1
      , (Product2_1_index_acc_sdt[0])});
  assign Accum2_mux_134_nl = MUX_v_16_2_2(Accum2_mux_135_nl, Accum2_1_mux_7_nl, fsm_output[11]);
  assign nl_z_out_6 = Accum2_mux_133_nl + Accum2_mux_134_nl;
  assign z_out_6 = nl_z_out_6[15:0];

  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_4_2;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [3:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    MUX1HOT_v_16_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_5_2;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [4:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    MUX1HOT_v_7_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_128_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [15:0] input_56;
    input [15:0] input_57;
    input [15:0] input_58;
    input [15:0] input_59;
    input [15:0] input_60;
    input [15:0] input_61;
    input [15:0] input_62;
    input [15:0] input_63;
    input [15:0] input_64;
    input [15:0] input_65;
    input [15:0] input_66;
    input [15:0] input_67;
    input [15:0] input_68;
    input [15:0] input_69;
    input [15:0] input_70;
    input [15:0] input_71;
    input [15:0] input_72;
    input [15:0] input_73;
    input [15:0] input_74;
    input [15:0] input_75;
    input [15:0] input_76;
    input [15:0] input_77;
    input [15:0] input_78;
    input [15:0] input_79;
    input [15:0] input_80;
    input [15:0] input_81;
    input [15:0] input_82;
    input [15:0] input_83;
    input [15:0] input_84;
    input [15:0] input_85;
    input [15:0] input_86;
    input [15:0] input_87;
    input [15:0] input_88;
    input [15:0] input_89;
    input [15:0] input_90;
    input [15:0] input_91;
    input [15:0] input_92;
    input [15:0] input_93;
    input [15:0] input_94;
    input [15:0] input_95;
    input [15:0] input_96;
    input [15:0] input_97;
    input [15:0] input_98;
    input [15:0] input_99;
    input [15:0] input_100;
    input [15:0] input_101;
    input [15:0] input_102;
    input [15:0] input_103;
    input [15:0] input_104;
    input [15:0] input_105;
    input [15:0] input_106;
    input [15:0] input_107;
    input [15:0] input_108;
    input [15:0] input_109;
    input [15:0] input_110;
    input [15:0] input_111;
    input [15:0] input_112;
    input [15:0] input_113;
    input [15:0] input_114;
    input [15:0] input_115;
    input [15:0] input_116;
    input [15:0] input_117;
    input [15:0] input_118;
    input [15:0] input_119;
    input [15:0] input_120;
    input [15:0] input_121;
    input [15:0] input_122;
    input [15:0] input_123;
    input [15:0] input_124;
    input [15:0] input_125;
    input [15:0] input_126;
    input [15:0] input_127;
    input [6:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      7'b1111101 : begin
        result = input_125;
      end
      7'b1111110 : begin
        result = input_126;
      end
      default : begin
        result = input_127;
      end
    endcase
    MUX_v_16_128_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_14_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [3:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      default : begin
        result = input_13;
      end
    endcase
    MUX_v_16_14_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_1792_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [15:0] input_56;
    input [15:0] input_57;
    input [15:0] input_58;
    input [15:0] input_59;
    input [15:0] input_60;
    input [15:0] input_61;
    input [15:0] input_62;
    input [15:0] input_63;
    input [15:0] input_64;
    input [15:0] input_65;
    input [15:0] input_66;
    input [15:0] input_67;
    input [15:0] input_68;
    input [15:0] input_69;
    input [15:0] input_70;
    input [15:0] input_71;
    input [15:0] input_72;
    input [15:0] input_73;
    input [15:0] input_74;
    input [15:0] input_75;
    input [15:0] input_76;
    input [15:0] input_77;
    input [15:0] input_78;
    input [15:0] input_79;
    input [15:0] input_80;
    input [15:0] input_81;
    input [15:0] input_82;
    input [15:0] input_83;
    input [15:0] input_84;
    input [15:0] input_85;
    input [15:0] input_86;
    input [15:0] input_87;
    input [15:0] input_88;
    input [15:0] input_89;
    input [15:0] input_90;
    input [15:0] input_91;
    input [15:0] input_92;
    input [15:0] input_93;
    input [15:0] input_94;
    input [15:0] input_95;
    input [15:0] input_96;
    input [15:0] input_97;
    input [15:0] input_98;
    input [15:0] input_99;
    input [15:0] input_100;
    input [15:0] input_101;
    input [15:0] input_102;
    input [15:0] input_103;
    input [15:0] input_104;
    input [15:0] input_105;
    input [15:0] input_106;
    input [15:0] input_107;
    input [15:0] input_108;
    input [15:0] input_109;
    input [15:0] input_110;
    input [15:0] input_111;
    input [15:0] input_112;
    input [15:0] input_113;
    input [15:0] input_114;
    input [15:0] input_115;
    input [15:0] input_116;
    input [15:0] input_117;
    input [15:0] input_118;
    input [15:0] input_119;
    input [15:0] input_120;
    input [15:0] input_121;
    input [15:0] input_122;
    input [15:0] input_123;
    input [15:0] input_124;
    input [15:0] input_125;
    input [15:0] input_126;
    input [15:0] input_127;
    input [15:0] input_128;
    input [15:0] input_129;
    input [15:0] input_130;
    input [15:0] input_131;
    input [15:0] input_132;
    input [15:0] input_133;
    input [15:0] input_134;
    input [15:0] input_135;
    input [15:0] input_136;
    input [15:0] input_137;
    input [15:0] input_138;
    input [15:0] input_139;
    input [15:0] input_140;
    input [15:0] input_141;
    input [15:0] input_142;
    input [15:0] input_143;
    input [15:0] input_144;
    input [15:0] input_145;
    input [15:0] input_146;
    input [15:0] input_147;
    input [15:0] input_148;
    input [15:0] input_149;
    input [15:0] input_150;
    input [15:0] input_151;
    input [15:0] input_152;
    input [15:0] input_153;
    input [15:0] input_154;
    input [15:0] input_155;
    input [15:0] input_156;
    input [15:0] input_157;
    input [15:0] input_158;
    input [15:0] input_159;
    input [15:0] input_160;
    input [15:0] input_161;
    input [15:0] input_162;
    input [15:0] input_163;
    input [15:0] input_164;
    input [15:0] input_165;
    input [15:0] input_166;
    input [15:0] input_167;
    input [15:0] input_168;
    input [15:0] input_169;
    input [15:0] input_170;
    input [15:0] input_171;
    input [15:0] input_172;
    input [15:0] input_173;
    input [15:0] input_174;
    input [15:0] input_175;
    input [15:0] input_176;
    input [15:0] input_177;
    input [15:0] input_178;
    input [15:0] input_179;
    input [15:0] input_180;
    input [15:0] input_181;
    input [15:0] input_182;
    input [15:0] input_183;
    input [15:0] input_184;
    input [15:0] input_185;
    input [15:0] input_186;
    input [15:0] input_187;
    input [15:0] input_188;
    input [15:0] input_189;
    input [15:0] input_190;
    input [15:0] input_191;
    input [15:0] input_192;
    input [15:0] input_193;
    input [15:0] input_194;
    input [15:0] input_195;
    input [15:0] input_196;
    input [15:0] input_197;
    input [15:0] input_198;
    input [15:0] input_199;
    input [15:0] input_200;
    input [15:0] input_201;
    input [15:0] input_202;
    input [15:0] input_203;
    input [15:0] input_204;
    input [15:0] input_205;
    input [15:0] input_206;
    input [15:0] input_207;
    input [15:0] input_208;
    input [15:0] input_209;
    input [15:0] input_210;
    input [15:0] input_211;
    input [15:0] input_212;
    input [15:0] input_213;
    input [15:0] input_214;
    input [15:0] input_215;
    input [15:0] input_216;
    input [15:0] input_217;
    input [15:0] input_218;
    input [15:0] input_219;
    input [15:0] input_220;
    input [15:0] input_221;
    input [15:0] input_222;
    input [15:0] input_223;
    input [15:0] input_224;
    input [15:0] input_225;
    input [15:0] input_226;
    input [15:0] input_227;
    input [15:0] input_228;
    input [15:0] input_229;
    input [15:0] input_230;
    input [15:0] input_231;
    input [15:0] input_232;
    input [15:0] input_233;
    input [15:0] input_234;
    input [15:0] input_235;
    input [15:0] input_236;
    input [15:0] input_237;
    input [15:0] input_238;
    input [15:0] input_239;
    input [15:0] input_240;
    input [15:0] input_241;
    input [15:0] input_242;
    input [15:0] input_243;
    input [15:0] input_244;
    input [15:0] input_245;
    input [15:0] input_246;
    input [15:0] input_247;
    input [15:0] input_248;
    input [15:0] input_249;
    input [15:0] input_250;
    input [15:0] input_251;
    input [15:0] input_252;
    input [15:0] input_253;
    input [15:0] input_254;
    input [15:0] input_255;
    input [15:0] input_256;
    input [15:0] input_257;
    input [15:0] input_258;
    input [15:0] input_259;
    input [15:0] input_260;
    input [15:0] input_261;
    input [15:0] input_262;
    input [15:0] input_263;
    input [15:0] input_264;
    input [15:0] input_265;
    input [15:0] input_266;
    input [15:0] input_267;
    input [15:0] input_268;
    input [15:0] input_269;
    input [15:0] input_270;
    input [15:0] input_271;
    input [15:0] input_272;
    input [15:0] input_273;
    input [15:0] input_274;
    input [15:0] input_275;
    input [15:0] input_276;
    input [15:0] input_277;
    input [15:0] input_278;
    input [15:0] input_279;
    input [15:0] input_280;
    input [15:0] input_281;
    input [15:0] input_282;
    input [15:0] input_283;
    input [15:0] input_284;
    input [15:0] input_285;
    input [15:0] input_286;
    input [15:0] input_287;
    input [15:0] input_288;
    input [15:0] input_289;
    input [15:0] input_290;
    input [15:0] input_291;
    input [15:0] input_292;
    input [15:0] input_293;
    input [15:0] input_294;
    input [15:0] input_295;
    input [15:0] input_296;
    input [15:0] input_297;
    input [15:0] input_298;
    input [15:0] input_299;
    input [15:0] input_300;
    input [15:0] input_301;
    input [15:0] input_302;
    input [15:0] input_303;
    input [15:0] input_304;
    input [15:0] input_305;
    input [15:0] input_306;
    input [15:0] input_307;
    input [15:0] input_308;
    input [15:0] input_309;
    input [15:0] input_310;
    input [15:0] input_311;
    input [15:0] input_312;
    input [15:0] input_313;
    input [15:0] input_314;
    input [15:0] input_315;
    input [15:0] input_316;
    input [15:0] input_317;
    input [15:0] input_318;
    input [15:0] input_319;
    input [15:0] input_320;
    input [15:0] input_321;
    input [15:0] input_322;
    input [15:0] input_323;
    input [15:0] input_324;
    input [15:0] input_325;
    input [15:0] input_326;
    input [15:0] input_327;
    input [15:0] input_328;
    input [15:0] input_329;
    input [15:0] input_330;
    input [15:0] input_331;
    input [15:0] input_332;
    input [15:0] input_333;
    input [15:0] input_334;
    input [15:0] input_335;
    input [15:0] input_336;
    input [15:0] input_337;
    input [15:0] input_338;
    input [15:0] input_339;
    input [15:0] input_340;
    input [15:0] input_341;
    input [15:0] input_342;
    input [15:0] input_343;
    input [15:0] input_344;
    input [15:0] input_345;
    input [15:0] input_346;
    input [15:0] input_347;
    input [15:0] input_348;
    input [15:0] input_349;
    input [15:0] input_350;
    input [15:0] input_351;
    input [15:0] input_352;
    input [15:0] input_353;
    input [15:0] input_354;
    input [15:0] input_355;
    input [15:0] input_356;
    input [15:0] input_357;
    input [15:0] input_358;
    input [15:0] input_359;
    input [15:0] input_360;
    input [15:0] input_361;
    input [15:0] input_362;
    input [15:0] input_363;
    input [15:0] input_364;
    input [15:0] input_365;
    input [15:0] input_366;
    input [15:0] input_367;
    input [15:0] input_368;
    input [15:0] input_369;
    input [15:0] input_370;
    input [15:0] input_371;
    input [15:0] input_372;
    input [15:0] input_373;
    input [15:0] input_374;
    input [15:0] input_375;
    input [15:0] input_376;
    input [15:0] input_377;
    input [15:0] input_378;
    input [15:0] input_379;
    input [15:0] input_380;
    input [15:0] input_381;
    input [15:0] input_382;
    input [15:0] input_383;
    input [15:0] input_384;
    input [15:0] input_385;
    input [15:0] input_386;
    input [15:0] input_387;
    input [15:0] input_388;
    input [15:0] input_389;
    input [15:0] input_390;
    input [15:0] input_391;
    input [15:0] input_392;
    input [15:0] input_393;
    input [15:0] input_394;
    input [15:0] input_395;
    input [15:0] input_396;
    input [15:0] input_397;
    input [15:0] input_398;
    input [15:0] input_399;
    input [15:0] input_400;
    input [15:0] input_401;
    input [15:0] input_402;
    input [15:0] input_403;
    input [15:0] input_404;
    input [15:0] input_405;
    input [15:0] input_406;
    input [15:0] input_407;
    input [15:0] input_408;
    input [15:0] input_409;
    input [15:0] input_410;
    input [15:0] input_411;
    input [15:0] input_412;
    input [15:0] input_413;
    input [15:0] input_414;
    input [15:0] input_415;
    input [15:0] input_416;
    input [15:0] input_417;
    input [15:0] input_418;
    input [15:0] input_419;
    input [15:0] input_420;
    input [15:0] input_421;
    input [15:0] input_422;
    input [15:0] input_423;
    input [15:0] input_424;
    input [15:0] input_425;
    input [15:0] input_426;
    input [15:0] input_427;
    input [15:0] input_428;
    input [15:0] input_429;
    input [15:0] input_430;
    input [15:0] input_431;
    input [15:0] input_432;
    input [15:0] input_433;
    input [15:0] input_434;
    input [15:0] input_435;
    input [15:0] input_436;
    input [15:0] input_437;
    input [15:0] input_438;
    input [15:0] input_439;
    input [15:0] input_440;
    input [15:0] input_441;
    input [15:0] input_442;
    input [15:0] input_443;
    input [15:0] input_444;
    input [15:0] input_445;
    input [15:0] input_446;
    input [15:0] input_447;
    input [15:0] input_448;
    input [15:0] input_449;
    input [15:0] input_450;
    input [15:0] input_451;
    input [15:0] input_452;
    input [15:0] input_453;
    input [15:0] input_454;
    input [15:0] input_455;
    input [15:0] input_456;
    input [15:0] input_457;
    input [15:0] input_458;
    input [15:0] input_459;
    input [15:0] input_460;
    input [15:0] input_461;
    input [15:0] input_462;
    input [15:0] input_463;
    input [15:0] input_464;
    input [15:0] input_465;
    input [15:0] input_466;
    input [15:0] input_467;
    input [15:0] input_468;
    input [15:0] input_469;
    input [15:0] input_470;
    input [15:0] input_471;
    input [15:0] input_472;
    input [15:0] input_473;
    input [15:0] input_474;
    input [15:0] input_475;
    input [15:0] input_476;
    input [15:0] input_477;
    input [15:0] input_478;
    input [15:0] input_479;
    input [15:0] input_480;
    input [15:0] input_481;
    input [15:0] input_482;
    input [15:0] input_483;
    input [15:0] input_484;
    input [15:0] input_485;
    input [15:0] input_486;
    input [15:0] input_487;
    input [15:0] input_488;
    input [15:0] input_489;
    input [15:0] input_490;
    input [15:0] input_491;
    input [15:0] input_492;
    input [15:0] input_493;
    input [15:0] input_494;
    input [15:0] input_495;
    input [15:0] input_496;
    input [15:0] input_497;
    input [15:0] input_498;
    input [15:0] input_499;
    input [15:0] input_500;
    input [15:0] input_501;
    input [15:0] input_502;
    input [15:0] input_503;
    input [15:0] input_504;
    input [15:0] input_505;
    input [15:0] input_506;
    input [15:0] input_507;
    input [15:0] input_508;
    input [15:0] input_509;
    input [15:0] input_510;
    input [15:0] input_511;
    input [15:0] input_512;
    input [15:0] input_513;
    input [15:0] input_514;
    input [15:0] input_515;
    input [15:0] input_516;
    input [15:0] input_517;
    input [15:0] input_518;
    input [15:0] input_519;
    input [15:0] input_520;
    input [15:0] input_521;
    input [15:0] input_522;
    input [15:0] input_523;
    input [15:0] input_524;
    input [15:0] input_525;
    input [15:0] input_526;
    input [15:0] input_527;
    input [15:0] input_528;
    input [15:0] input_529;
    input [15:0] input_530;
    input [15:0] input_531;
    input [15:0] input_532;
    input [15:0] input_533;
    input [15:0] input_534;
    input [15:0] input_535;
    input [15:0] input_536;
    input [15:0] input_537;
    input [15:0] input_538;
    input [15:0] input_539;
    input [15:0] input_540;
    input [15:0] input_541;
    input [15:0] input_542;
    input [15:0] input_543;
    input [15:0] input_544;
    input [15:0] input_545;
    input [15:0] input_546;
    input [15:0] input_547;
    input [15:0] input_548;
    input [15:0] input_549;
    input [15:0] input_550;
    input [15:0] input_551;
    input [15:0] input_552;
    input [15:0] input_553;
    input [15:0] input_554;
    input [15:0] input_555;
    input [15:0] input_556;
    input [15:0] input_557;
    input [15:0] input_558;
    input [15:0] input_559;
    input [15:0] input_560;
    input [15:0] input_561;
    input [15:0] input_562;
    input [15:0] input_563;
    input [15:0] input_564;
    input [15:0] input_565;
    input [15:0] input_566;
    input [15:0] input_567;
    input [15:0] input_568;
    input [15:0] input_569;
    input [15:0] input_570;
    input [15:0] input_571;
    input [15:0] input_572;
    input [15:0] input_573;
    input [15:0] input_574;
    input [15:0] input_575;
    input [15:0] input_576;
    input [15:0] input_577;
    input [15:0] input_578;
    input [15:0] input_579;
    input [15:0] input_580;
    input [15:0] input_581;
    input [15:0] input_582;
    input [15:0] input_583;
    input [15:0] input_584;
    input [15:0] input_585;
    input [15:0] input_586;
    input [15:0] input_587;
    input [15:0] input_588;
    input [15:0] input_589;
    input [15:0] input_590;
    input [15:0] input_591;
    input [15:0] input_592;
    input [15:0] input_593;
    input [15:0] input_594;
    input [15:0] input_595;
    input [15:0] input_596;
    input [15:0] input_597;
    input [15:0] input_598;
    input [15:0] input_599;
    input [15:0] input_600;
    input [15:0] input_601;
    input [15:0] input_602;
    input [15:0] input_603;
    input [15:0] input_604;
    input [15:0] input_605;
    input [15:0] input_606;
    input [15:0] input_607;
    input [15:0] input_608;
    input [15:0] input_609;
    input [15:0] input_610;
    input [15:0] input_611;
    input [15:0] input_612;
    input [15:0] input_613;
    input [15:0] input_614;
    input [15:0] input_615;
    input [15:0] input_616;
    input [15:0] input_617;
    input [15:0] input_618;
    input [15:0] input_619;
    input [15:0] input_620;
    input [15:0] input_621;
    input [15:0] input_622;
    input [15:0] input_623;
    input [15:0] input_624;
    input [15:0] input_625;
    input [15:0] input_626;
    input [15:0] input_627;
    input [15:0] input_628;
    input [15:0] input_629;
    input [15:0] input_630;
    input [15:0] input_631;
    input [15:0] input_632;
    input [15:0] input_633;
    input [15:0] input_634;
    input [15:0] input_635;
    input [15:0] input_636;
    input [15:0] input_637;
    input [15:0] input_638;
    input [15:0] input_639;
    input [15:0] input_640;
    input [15:0] input_641;
    input [15:0] input_642;
    input [15:0] input_643;
    input [15:0] input_644;
    input [15:0] input_645;
    input [15:0] input_646;
    input [15:0] input_647;
    input [15:0] input_648;
    input [15:0] input_649;
    input [15:0] input_650;
    input [15:0] input_651;
    input [15:0] input_652;
    input [15:0] input_653;
    input [15:0] input_654;
    input [15:0] input_655;
    input [15:0] input_656;
    input [15:0] input_657;
    input [15:0] input_658;
    input [15:0] input_659;
    input [15:0] input_660;
    input [15:0] input_661;
    input [15:0] input_662;
    input [15:0] input_663;
    input [15:0] input_664;
    input [15:0] input_665;
    input [15:0] input_666;
    input [15:0] input_667;
    input [15:0] input_668;
    input [15:0] input_669;
    input [15:0] input_670;
    input [15:0] input_671;
    input [15:0] input_672;
    input [15:0] input_673;
    input [15:0] input_674;
    input [15:0] input_675;
    input [15:0] input_676;
    input [15:0] input_677;
    input [15:0] input_678;
    input [15:0] input_679;
    input [15:0] input_680;
    input [15:0] input_681;
    input [15:0] input_682;
    input [15:0] input_683;
    input [15:0] input_684;
    input [15:0] input_685;
    input [15:0] input_686;
    input [15:0] input_687;
    input [15:0] input_688;
    input [15:0] input_689;
    input [15:0] input_690;
    input [15:0] input_691;
    input [15:0] input_692;
    input [15:0] input_693;
    input [15:0] input_694;
    input [15:0] input_695;
    input [15:0] input_696;
    input [15:0] input_697;
    input [15:0] input_698;
    input [15:0] input_699;
    input [15:0] input_700;
    input [15:0] input_701;
    input [15:0] input_702;
    input [15:0] input_703;
    input [15:0] input_704;
    input [15:0] input_705;
    input [15:0] input_706;
    input [15:0] input_707;
    input [15:0] input_708;
    input [15:0] input_709;
    input [15:0] input_710;
    input [15:0] input_711;
    input [15:0] input_712;
    input [15:0] input_713;
    input [15:0] input_714;
    input [15:0] input_715;
    input [15:0] input_716;
    input [15:0] input_717;
    input [15:0] input_718;
    input [15:0] input_719;
    input [15:0] input_720;
    input [15:0] input_721;
    input [15:0] input_722;
    input [15:0] input_723;
    input [15:0] input_724;
    input [15:0] input_725;
    input [15:0] input_726;
    input [15:0] input_727;
    input [15:0] input_728;
    input [15:0] input_729;
    input [15:0] input_730;
    input [15:0] input_731;
    input [15:0] input_732;
    input [15:0] input_733;
    input [15:0] input_734;
    input [15:0] input_735;
    input [15:0] input_736;
    input [15:0] input_737;
    input [15:0] input_738;
    input [15:0] input_739;
    input [15:0] input_740;
    input [15:0] input_741;
    input [15:0] input_742;
    input [15:0] input_743;
    input [15:0] input_744;
    input [15:0] input_745;
    input [15:0] input_746;
    input [15:0] input_747;
    input [15:0] input_748;
    input [15:0] input_749;
    input [15:0] input_750;
    input [15:0] input_751;
    input [15:0] input_752;
    input [15:0] input_753;
    input [15:0] input_754;
    input [15:0] input_755;
    input [15:0] input_756;
    input [15:0] input_757;
    input [15:0] input_758;
    input [15:0] input_759;
    input [15:0] input_760;
    input [15:0] input_761;
    input [15:0] input_762;
    input [15:0] input_763;
    input [15:0] input_764;
    input [15:0] input_765;
    input [15:0] input_766;
    input [15:0] input_767;
    input [15:0] input_768;
    input [15:0] input_769;
    input [15:0] input_770;
    input [15:0] input_771;
    input [15:0] input_772;
    input [15:0] input_773;
    input [15:0] input_774;
    input [15:0] input_775;
    input [15:0] input_776;
    input [15:0] input_777;
    input [15:0] input_778;
    input [15:0] input_779;
    input [15:0] input_780;
    input [15:0] input_781;
    input [15:0] input_782;
    input [15:0] input_783;
    input [15:0] input_784;
    input [15:0] input_785;
    input [15:0] input_786;
    input [15:0] input_787;
    input [15:0] input_788;
    input [15:0] input_789;
    input [15:0] input_790;
    input [15:0] input_791;
    input [15:0] input_792;
    input [15:0] input_793;
    input [15:0] input_794;
    input [15:0] input_795;
    input [15:0] input_796;
    input [15:0] input_797;
    input [15:0] input_798;
    input [15:0] input_799;
    input [15:0] input_800;
    input [15:0] input_801;
    input [15:0] input_802;
    input [15:0] input_803;
    input [15:0] input_804;
    input [15:0] input_805;
    input [15:0] input_806;
    input [15:0] input_807;
    input [15:0] input_808;
    input [15:0] input_809;
    input [15:0] input_810;
    input [15:0] input_811;
    input [15:0] input_812;
    input [15:0] input_813;
    input [15:0] input_814;
    input [15:0] input_815;
    input [15:0] input_816;
    input [15:0] input_817;
    input [15:0] input_818;
    input [15:0] input_819;
    input [15:0] input_820;
    input [15:0] input_821;
    input [15:0] input_822;
    input [15:0] input_823;
    input [15:0] input_824;
    input [15:0] input_825;
    input [15:0] input_826;
    input [15:0] input_827;
    input [15:0] input_828;
    input [15:0] input_829;
    input [15:0] input_830;
    input [15:0] input_831;
    input [15:0] input_832;
    input [15:0] input_833;
    input [15:0] input_834;
    input [15:0] input_835;
    input [15:0] input_836;
    input [15:0] input_837;
    input [15:0] input_838;
    input [15:0] input_839;
    input [15:0] input_840;
    input [15:0] input_841;
    input [15:0] input_842;
    input [15:0] input_843;
    input [15:0] input_844;
    input [15:0] input_845;
    input [15:0] input_846;
    input [15:0] input_847;
    input [15:0] input_848;
    input [15:0] input_849;
    input [15:0] input_850;
    input [15:0] input_851;
    input [15:0] input_852;
    input [15:0] input_853;
    input [15:0] input_854;
    input [15:0] input_855;
    input [15:0] input_856;
    input [15:0] input_857;
    input [15:0] input_858;
    input [15:0] input_859;
    input [15:0] input_860;
    input [15:0] input_861;
    input [15:0] input_862;
    input [15:0] input_863;
    input [15:0] input_864;
    input [15:0] input_865;
    input [15:0] input_866;
    input [15:0] input_867;
    input [15:0] input_868;
    input [15:0] input_869;
    input [15:0] input_870;
    input [15:0] input_871;
    input [15:0] input_872;
    input [15:0] input_873;
    input [15:0] input_874;
    input [15:0] input_875;
    input [15:0] input_876;
    input [15:0] input_877;
    input [15:0] input_878;
    input [15:0] input_879;
    input [15:0] input_880;
    input [15:0] input_881;
    input [15:0] input_882;
    input [15:0] input_883;
    input [15:0] input_884;
    input [15:0] input_885;
    input [15:0] input_886;
    input [15:0] input_887;
    input [15:0] input_888;
    input [15:0] input_889;
    input [15:0] input_890;
    input [15:0] input_891;
    input [15:0] input_892;
    input [15:0] input_893;
    input [15:0] input_894;
    input [15:0] input_895;
    input [15:0] input_896;
    input [15:0] input_897;
    input [15:0] input_898;
    input [15:0] input_899;
    input [15:0] input_900;
    input [15:0] input_901;
    input [15:0] input_902;
    input [15:0] input_903;
    input [15:0] input_904;
    input [15:0] input_905;
    input [15:0] input_906;
    input [15:0] input_907;
    input [15:0] input_908;
    input [15:0] input_909;
    input [15:0] input_910;
    input [15:0] input_911;
    input [15:0] input_912;
    input [15:0] input_913;
    input [15:0] input_914;
    input [15:0] input_915;
    input [15:0] input_916;
    input [15:0] input_917;
    input [15:0] input_918;
    input [15:0] input_919;
    input [15:0] input_920;
    input [15:0] input_921;
    input [15:0] input_922;
    input [15:0] input_923;
    input [15:0] input_924;
    input [15:0] input_925;
    input [15:0] input_926;
    input [15:0] input_927;
    input [15:0] input_928;
    input [15:0] input_929;
    input [15:0] input_930;
    input [15:0] input_931;
    input [15:0] input_932;
    input [15:0] input_933;
    input [15:0] input_934;
    input [15:0] input_935;
    input [15:0] input_936;
    input [15:0] input_937;
    input [15:0] input_938;
    input [15:0] input_939;
    input [15:0] input_940;
    input [15:0] input_941;
    input [15:0] input_942;
    input [15:0] input_943;
    input [15:0] input_944;
    input [15:0] input_945;
    input [15:0] input_946;
    input [15:0] input_947;
    input [15:0] input_948;
    input [15:0] input_949;
    input [15:0] input_950;
    input [15:0] input_951;
    input [15:0] input_952;
    input [15:0] input_953;
    input [15:0] input_954;
    input [15:0] input_955;
    input [15:0] input_956;
    input [15:0] input_957;
    input [15:0] input_958;
    input [15:0] input_959;
    input [15:0] input_960;
    input [15:0] input_961;
    input [15:0] input_962;
    input [15:0] input_963;
    input [15:0] input_964;
    input [15:0] input_965;
    input [15:0] input_966;
    input [15:0] input_967;
    input [15:0] input_968;
    input [15:0] input_969;
    input [15:0] input_970;
    input [15:0] input_971;
    input [15:0] input_972;
    input [15:0] input_973;
    input [15:0] input_974;
    input [15:0] input_975;
    input [15:0] input_976;
    input [15:0] input_977;
    input [15:0] input_978;
    input [15:0] input_979;
    input [15:0] input_980;
    input [15:0] input_981;
    input [15:0] input_982;
    input [15:0] input_983;
    input [15:0] input_984;
    input [15:0] input_985;
    input [15:0] input_986;
    input [15:0] input_987;
    input [15:0] input_988;
    input [15:0] input_989;
    input [15:0] input_990;
    input [15:0] input_991;
    input [15:0] input_992;
    input [15:0] input_993;
    input [15:0] input_994;
    input [15:0] input_995;
    input [15:0] input_996;
    input [15:0] input_997;
    input [15:0] input_998;
    input [15:0] input_999;
    input [15:0] input_1000;
    input [15:0] input_1001;
    input [15:0] input_1002;
    input [15:0] input_1003;
    input [15:0] input_1004;
    input [15:0] input_1005;
    input [15:0] input_1006;
    input [15:0] input_1007;
    input [15:0] input_1008;
    input [15:0] input_1009;
    input [15:0] input_1010;
    input [15:0] input_1011;
    input [15:0] input_1012;
    input [15:0] input_1013;
    input [15:0] input_1014;
    input [15:0] input_1015;
    input [15:0] input_1016;
    input [15:0] input_1017;
    input [15:0] input_1018;
    input [15:0] input_1019;
    input [15:0] input_1020;
    input [15:0] input_1021;
    input [15:0] input_1022;
    input [15:0] input_1023;
    input [15:0] input_1024;
    input [15:0] input_1025;
    input [15:0] input_1026;
    input [15:0] input_1027;
    input [15:0] input_1028;
    input [15:0] input_1029;
    input [15:0] input_1030;
    input [15:0] input_1031;
    input [15:0] input_1032;
    input [15:0] input_1033;
    input [15:0] input_1034;
    input [15:0] input_1035;
    input [15:0] input_1036;
    input [15:0] input_1037;
    input [15:0] input_1038;
    input [15:0] input_1039;
    input [15:0] input_1040;
    input [15:0] input_1041;
    input [15:0] input_1042;
    input [15:0] input_1043;
    input [15:0] input_1044;
    input [15:0] input_1045;
    input [15:0] input_1046;
    input [15:0] input_1047;
    input [15:0] input_1048;
    input [15:0] input_1049;
    input [15:0] input_1050;
    input [15:0] input_1051;
    input [15:0] input_1052;
    input [15:0] input_1053;
    input [15:0] input_1054;
    input [15:0] input_1055;
    input [15:0] input_1056;
    input [15:0] input_1057;
    input [15:0] input_1058;
    input [15:0] input_1059;
    input [15:0] input_1060;
    input [15:0] input_1061;
    input [15:0] input_1062;
    input [15:0] input_1063;
    input [15:0] input_1064;
    input [15:0] input_1065;
    input [15:0] input_1066;
    input [15:0] input_1067;
    input [15:0] input_1068;
    input [15:0] input_1069;
    input [15:0] input_1070;
    input [15:0] input_1071;
    input [15:0] input_1072;
    input [15:0] input_1073;
    input [15:0] input_1074;
    input [15:0] input_1075;
    input [15:0] input_1076;
    input [15:0] input_1077;
    input [15:0] input_1078;
    input [15:0] input_1079;
    input [15:0] input_1080;
    input [15:0] input_1081;
    input [15:0] input_1082;
    input [15:0] input_1083;
    input [15:0] input_1084;
    input [15:0] input_1085;
    input [15:0] input_1086;
    input [15:0] input_1087;
    input [15:0] input_1088;
    input [15:0] input_1089;
    input [15:0] input_1090;
    input [15:0] input_1091;
    input [15:0] input_1092;
    input [15:0] input_1093;
    input [15:0] input_1094;
    input [15:0] input_1095;
    input [15:0] input_1096;
    input [15:0] input_1097;
    input [15:0] input_1098;
    input [15:0] input_1099;
    input [15:0] input_1100;
    input [15:0] input_1101;
    input [15:0] input_1102;
    input [15:0] input_1103;
    input [15:0] input_1104;
    input [15:0] input_1105;
    input [15:0] input_1106;
    input [15:0] input_1107;
    input [15:0] input_1108;
    input [15:0] input_1109;
    input [15:0] input_1110;
    input [15:0] input_1111;
    input [15:0] input_1112;
    input [15:0] input_1113;
    input [15:0] input_1114;
    input [15:0] input_1115;
    input [15:0] input_1116;
    input [15:0] input_1117;
    input [15:0] input_1118;
    input [15:0] input_1119;
    input [15:0] input_1120;
    input [15:0] input_1121;
    input [15:0] input_1122;
    input [15:0] input_1123;
    input [15:0] input_1124;
    input [15:0] input_1125;
    input [15:0] input_1126;
    input [15:0] input_1127;
    input [15:0] input_1128;
    input [15:0] input_1129;
    input [15:0] input_1130;
    input [15:0] input_1131;
    input [15:0] input_1132;
    input [15:0] input_1133;
    input [15:0] input_1134;
    input [15:0] input_1135;
    input [15:0] input_1136;
    input [15:0] input_1137;
    input [15:0] input_1138;
    input [15:0] input_1139;
    input [15:0] input_1140;
    input [15:0] input_1141;
    input [15:0] input_1142;
    input [15:0] input_1143;
    input [15:0] input_1144;
    input [15:0] input_1145;
    input [15:0] input_1146;
    input [15:0] input_1147;
    input [15:0] input_1148;
    input [15:0] input_1149;
    input [15:0] input_1150;
    input [15:0] input_1151;
    input [15:0] input_1152;
    input [15:0] input_1153;
    input [15:0] input_1154;
    input [15:0] input_1155;
    input [15:0] input_1156;
    input [15:0] input_1157;
    input [15:0] input_1158;
    input [15:0] input_1159;
    input [15:0] input_1160;
    input [15:0] input_1161;
    input [15:0] input_1162;
    input [15:0] input_1163;
    input [15:0] input_1164;
    input [15:0] input_1165;
    input [15:0] input_1166;
    input [15:0] input_1167;
    input [15:0] input_1168;
    input [15:0] input_1169;
    input [15:0] input_1170;
    input [15:0] input_1171;
    input [15:0] input_1172;
    input [15:0] input_1173;
    input [15:0] input_1174;
    input [15:0] input_1175;
    input [15:0] input_1176;
    input [15:0] input_1177;
    input [15:0] input_1178;
    input [15:0] input_1179;
    input [15:0] input_1180;
    input [15:0] input_1181;
    input [15:0] input_1182;
    input [15:0] input_1183;
    input [15:0] input_1184;
    input [15:0] input_1185;
    input [15:0] input_1186;
    input [15:0] input_1187;
    input [15:0] input_1188;
    input [15:0] input_1189;
    input [15:0] input_1190;
    input [15:0] input_1191;
    input [15:0] input_1192;
    input [15:0] input_1193;
    input [15:0] input_1194;
    input [15:0] input_1195;
    input [15:0] input_1196;
    input [15:0] input_1197;
    input [15:0] input_1198;
    input [15:0] input_1199;
    input [15:0] input_1200;
    input [15:0] input_1201;
    input [15:0] input_1202;
    input [15:0] input_1203;
    input [15:0] input_1204;
    input [15:0] input_1205;
    input [15:0] input_1206;
    input [15:0] input_1207;
    input [15:0] input_1208;
    input [15:0] input_1209;
    input [15:0] input_1210;
    input [15:0] input_1211;
    input [15:0] input_1212;
    input [15:0] input_1213;
    input [15:0] input_1214;
    input [15:0] input_1215;
    input [15:0] input_1216;
    input [15:0] input_1217;
    input [15:0] input_1218;
    input [15:0] input_1219;
    input [15:0] input_1220;
    input [15:0] input_1221;
    input [15:0] input_1222;
    input [15:0] input_1223;
    input [15:0] input_1224;
    input [15:0] input_1225;
    input [15:0] input_1226;
    input [15:0] input_1227;
    input [15:0] input_1228;
    input [15:0] input_1229;
    input [15:0] input_1230;
    input [15:0] input_1231;
    input [15:0] input_1232;
    input [15:0] input_1233;
    input [15:0] input_1234;
    input [15:0] input_1235;
    input [15:0] input_1236;
    input [15:0] input_1237;
    input [15:0] input_1238;
    input [15:0] input_1239;
    input [15:0] input_1240;
    input [15:0] input_1241;
    input [15:0] input_1242;
    input [15:0] input_1243;
    input [15:0] input_1244;
    input [15:0] input_1245;
    input [15:0] input_1246;
    input [15:0] input_1247;
    input [15:0] input_1248;
    input [15:0] input_1249;
    input [15:0] input_1250;
    input [15:0] input_1251;
    input [15:0] input_1252;
    input [15:0] input_1253;
    input [15:0] input_1254;
    input [15:0] input_1255;
    input [15:0] input_1256;
    input [15:0] input_1257;
    input [15:0] input_1258;
    input [15:0] input_1259;
    input [15:0] input_1260;
    input [15:0] input_1261;
    input [15:0] input_1262;
    input [15:0] input_1263;
    input [15:0] input_1264;
    input [15:0] input_1265;
    input [15:0] input_1266;
    input [15:0] input_1267;
    input [15:0] input_1268;
    input [15:0] input_1269;
    input [15:0] input_1270;
    input [15:0] input_1271;
    input [15:0] input_1272;
    input [15:0] input_1273;
    input [15:0] input_1274;
    input [15:0] input_1275;
    input [15:0] input_1276;
    input [15:0] input_1277;
    input [15:0] input_1278;
    input [15:0] input_1279;
    input [15:0] input_1280;
    input [15:0] input_1281;
    input [15:0] input_1282;
    input [15:0] input_1283;
    input [15:0] input_1284;
    input [15:0] input_1285;
    input [15:0] input_1286;
    input [15:0] input_1287;
    input [15:0] input_1288;
    input [15:0] input_1289;
    input [15:0] input_1290;
    input [15:0] input_1291;
    input [15:0] input_1292;
    input [15:0] input_1293;
    input [15:0] input_1294;
    input [15:0] input_1295;
    input [15:0] input_1296;
    input [15:0] input_1297;
    input [15:0] input_1298;
    input [15:0] input_1299;
    input [15:0] input_1300;
    input [15:0] input_1301;
    input [15:0] input_1302;
    input [15:0] input_1303;
    input [15:0] input_1304;
    input [15:0] input_1305;
    input [15:0] input_1306;
    input [15:0] input_1307;
    input [15:0] input_1308;
    input [15:0] input_1309;
    input [15:0] input_1310;
    input [15:0] input_1311;
    input [15:0] input_1312;
    input [15:0] input_1313;
    input [15:0] input_1314;
    input [15:0] input_1315;
    input [15:0] input_1316;
    input [15:0] input_1317;
    input [15:0] input_1318;
    input [15:0] input_1319;
    input [15:0] input_1320;
    input [15:0] input_1321;
    input [15:0] input_1322;
    input [15:0] input_1323;
    input [15:0] input_1324;
    input [15:0] input_1325;
    input [15:0] input_1326;
    input [15:0] input_1327;
    input [15:0] input_1328;
    input [15:0] input_1329;
    input [15:0] input_1330;
    input [15:0] input_1331;
    input [15:0] input_1332;
    input [15:0] input_1333;
    input [15:0] input_1334;
    input [15:0] input_1335;
    input [15:0] input_1336;
    input [15:0] input_1337;
    input [15:0] input_1338;
    input [15:0] input_1339;
    input [15:0] input_1340;
    input [15:0] input_1341;
    input [15:0] input_1342;
    input [15:0] input_1343;
    input [15:0] input_1344;
    input [15:0] input_1345;
    input [15:0] input_1346;
    input [15:0] input_1347;
    input [15:0] input_1348;
    input [15:0] input_1349;
    input [15:0] input_1350;
    input [15:0] input_1351;
    input [15:0] input_1352;
    input [15:0] input_1353;
    input [15:0] input_1354;
    input [15:0] input_1355;
    input [15:0] input_1356;
    input [15:0] input_1357;
    input [15:0] input_1358;
    input [15:0] input_1359;
    input [15:0] input_1360;
    input [15:0] input_1361;
    input [15:0] input_1362;
    input [15:0] input_1363;
    input [15:0] input_1364;
    input [15:0] input_1365;
    input [15:0] input_1366;
    input [15:0] input_1367;
    input [15:0] input_1368;
    input [15:0] input_1369;
    input [15:0] input_1370;
    input [15:0] input_1371;
    input [15:0] input_1372;
    input [15:0] input_1373;
    input [15:0] input_1374;
    input [15:0] input_1375;
    input [15:0] input_1376;
    input [15:0] input_1377;
    input [15:0] input_1378;
    input [15:0] input_1379;
    input [15:0] input_1380;
    input [15:0] input_1381;
    input [15:0] input_1382;
    input [15:0] input_1383;
    input [15:0] input_1384;
    input [15:0] input_1385;
    input [15:0] input_1386;
    input [15:0] input_1387;
    input [15:0] input_1388;
    input [15:0] input_1389;
    input [15:0] input_1390;
    input [15:0] input_1391;
    input [15:0] input_1392;
    input [15:0] input_1393;
    input [15:0] input_1394;
    input [15:0] input_1395;
    input [15:0] input_1396;
    input [15:0] input_1397;
    input [15:0] input_1398;
    input [15:0] input_1399;
    input [15:0] input_1400;
    input [15:0] input_1401;
    input [15:0] input_1402;
    input [15:0] input_1403;
    input [15:0] input_1404;
    input [15:0] input_1405;
    input [15:0] input_1406;
    input [15:0] input_1407;
    input [15:0] input_1408;
    input [15:0] input_1409;
    input [15:0] input_1410;
    input [15:0] input_1411;
    input [15:0] input_1412;
    input [15:0] input_1413;
    input [15:0] input_1414;
    input [15:0] input_1415;
    input [15:0] input_1416;
    input [15:0] input_1417;
    input [15:0] input_1418;
    input [15:0] input_1419;
    input [15:0] input_1420;
    input [15:0] input_1421;
    input [15:0] input_1422;
    input [15:0] input_1423;
    input [15:0] input_1424;
    input [15:0] input_1425;
    input [15:0] input_1426;
    input [15:0] input_1427;
    input [15:0] input_1428;
    input [15:0] input_1429;
    input [15:0] input_1430;
    input [15:0] input_1431;
    input [15:0] input_1432;
    input [15:0] input_1433;
    input [15:0] input_1434;
    input [15:0] input_1435;
    input [15:0] input_1436;
    input [15:0] input_1437;
    input [15:0] input_1438;
    input [15:0] input_1439;
    input [15:0] input_1440;
    input [15:0] input_1441;
    input [15:0] input_1442;
    input [15:0] input_1443;
    input [15:0] input_1444;
    input [15:0] input_1445;
    input [15:0] input_1446;
    input [15:0] input_1447;
    input [15:0] input_1448;
    input [15:0] input_1449;
    input [15:0] input_1450;
    input [15:0] input_1451;
    input [15:0] input_1452;
    input [15:0] input_1453;
    input [15:0] input_1454;
    input [15:0] input_1455;
    input [15:0] input_1456;
    input [15:0] input_1457;
    input [15:0] input_1458;
    input [15:0] input_1459;
    input [15:0] input_1460;
    input [15:0] input_1461;
    input [15:0] input_1462;
    input [15:0] input_1463;
    input [15:0] input_1464;
    input [15:0] input_1465;
    input [15:0] input_1466;
    input [15:0] input_1467;
    input [15:0] input_1468;
    input [15:0] input_1469;
    input [15:0] input_1470;
    input [15:0] input_1471;
    input [15:0] input_1472;
    input [15:0] input_1473;
    input [15:0] input_1474;
    input [15:0] input_1475;
    input [15:0] input_1476;
    input [15:0] input_1477;
    input [15:0] input_1478;
    input [15:0] input_1479;
    input [15:0] input_1480;
    input [15:0] input_1481;
    input [15:0] input_1482;
    input [15:0] input_1483;
    input [15:0] input_1484;
    input [15:0] input_1485;
    input [15:0] input_1486;
    input [15:0] input_1487;
    input [15:0] input_1488;
    input [15:0] input_1489;
    input [15:0] input_1490;
    input [15:0] input_1491;
    input [15:0] input_1492;
    input [15:0] input_1493;
    input [15:0] input_1494;
    input [15:0] input_1495;
    input [15:0] input_1496;
    input [15:0] input_1497;
    input [15:0] input_1498;
    input [15:0] input_1499;
    input [15:0] input_1500;
    input [15:0] input_1501;
    input [15:0] input_1502;
    input [15:0] input_1503;
    input [15:0] input_1504;
    input [15:0] input_1505;
    input [15:0] input_1506;
    input [15:0] input_1507;
    input [15:0] input_1508;
    input [15:0] input_1509;
    input [15:0] input_1510;
    input [15:0] input_1511;
    input [15:0] input_1512;
    input [15:0] input_1513;
    input [15:0] input_1514;
    input [15:0] input_1515;
    input [15:0] input_1516;
    input [15:0] input_1517;
    input [15:0] input_1518;
    input [15:0] input_1519;
    input [15:0] input_1520;
    input [15:0] input_1521;
    input [15:0] input_1522;
    input [15:0] input_1523;
    input [15:0] input_1524;
    input [15:0] input_1525;
    input [15:0] input_1526;
    input [15:0] input_1527;
    input [15:0] input_1528;
    input [15:0] input_1529;
    input [15:0] input_1530;
    input [15:0] input_1531;
    input [15:0] input_1532;
    input [15:0] input_1533;
    input [15:0] input_1534;
    input [15:0] input_1535;
    input [15:0] input_1536;
    input [15:0] input_1537;
    input [15:0] input_1538;
    input [15:0] input_1539;
    input [15:0] input_1540;
    input [15:0] input_1541;
    input [15:0] input_1542;
    input [15:0] input_1543;
    input [15:0] input_1544;
    input [15:0] input_1545;
    input [15:0] input_1546;
    input [15:0] input_1547;
    input [15:0] input_1548;
    input [15:0] input_1549;
    input [15:0] input_1550;
    input [15:0] input_1551;
    input [15:0] input_1552;
    input [15:0] input_1553;
    input [15:0] input_1554;
    input [15:0] input_1555;
    input [15:0] input_1556;
    input [15:0] input_1557;
    input [15:0] input_1558;
    input [15:0] input_1559;
    input [15:0] input_1560;
    input [15:0] input_1561;
    input [15:0] input_1562;
    input [15:0] input_1563;
    input [15:0] input_1564;
    input [15:0] input_1565;
    input [15:0] input_1566;
    input [15:0] input_1567;
    input [15:0] input_1568;
    input [15:0] input_1569;
    input [15:0] input_1570;
    input [15:0] input_1571;
    input [15:0] input_1572;
    input [15:0] input_1573;
    input [15:0] input_1574;
    input [15:0] input_1575;
    input [15:0] input_1576;
    input [15:0] input_1577;
    input [15:0] input_1578;
    input [15:0] input_1579;
    input [15:0] input_1580;
    input [15:0] input_1581;
    input [15:0] input_1582;
    input [15:0] input_1583;
    input [15:0] input_1584;
    input [15:0] input_1585;
    input [15:0] input_1586;
    input [15:0] input_1587;
    input [15:0] input_1588;
    input [15:0] input_1589;
    input [15:0] input_1590;
    input [15:0] input_1591;
    input [15:0] input_1592;
    input [15:0] input_1593;
    input [15:0] input_1594;
    input [15:0] input_1595;
    input [15:0] input_1596;
    input [15:0] input_1597;
    input [15:0] input_1598;
    input [15:0] input_1599;
    input [15:0] input_1600;
    input [15:0] input_1601;
    input [15:0] input_1602;
    input [15:0] input_1603;
    input [15:0] input_1604;
    input [15:0] input_1605;
    input [15:0] input_1606;
    input [15:0] input_1607;
    input [15:0] input_1608;
    input [15:0] input_1609;
    input [15:0] input_1610;
    input [15:0] input_1611;
    input [15:0] input_1612;
    input [15:0] input_1613;
    input [15:0] input_1614;
    input [15:0] input_1615;
    input [15:0] input_1616;
    input [15:0] input_1617;
    input [15:0] input_1618;
    input [15:0] input_1619;
    input [15:0] input_1620;
    input [15:0] input_1621;
    input [15:0] input_1622;
    input [15:0] input_1623;
    input [15:0] input_1624;
    input [15:0] input_1625;
    input [15:0] input_1626;
    input [15:0] input_1627;
    input [15:0] input_1628;
    input [15:0] input_1629;
    input [15:0] input_1630;
    input [15:0] input_1631;
    input [15:0] input_1632;
    input [15:0] input_1633;
    input [15:0] input_1634;
    input [15:0] input_1635;
    input [15:0] input_1636;
    input [15:0] input_1637;
    input [15:0] input_1638;
    input [15:0] input_1639;
    input [15:0] input_1640;
    input [15:0] input_1641;
    input [15:0] input_1642;
    input [15:0] input_1643;
    input [15:0] input_1644;
    input [15:0] input_1645;
    input [15:0] input_1646;
    input [15:0] input_1647;
    input [15:0] input_1648;
    input [15:0] input_1649;
    input [15:0] input_1650;
    input [15:0] input_1651;
    input [15:0] input_1652;
    input [15:0] input_1653;
    input [15:0] input_1654;
    input [15:0] input_1655;
    input [15:0] input_1656;
    input [15:0] input_1657;
    input [15:0] input_1658;
    input [15:0] input_1659;
    input [15:0] input_1660;
    input [15:0] input_1661;
    input [15:0] input_1662;
    input [15:0] input_1663;
    input [15:0] input_1664;
    input [15:0] input_1665;
    input [15:0] input_1666;
    input [15:0] input_1667;
    input [15:0] input_1668;
    input [15:0] input_1669;
    input [15:0] input_1670;
    input [15:0] input_1671;
    input [15:0] input_1672;
    input [15:0] input_1673;
    input [15:0] input_1674;
    input [15:0] input_1675;
    input [15:0] input_1676;
    input [15:0] input_1677;
    input [15:0] input_1678;
    input [15:0] input_1679;
    input [15:0] input_1680;
    input [15:0] input_1681;
    input [15:0] input_1682;
    input [15:0] input_1683;
    input [15:0] input_1684;
    input [15:0] input_1685;
    input [15:0] input_1686;
    input [15:0] input_1687;
    input [15:0] input_1688;
    input [15:0] input_1689;
    input [15:0] input_1690;
    input [15:0] input_1691;
    input [15:0] input_1692;
    input [15:0] input_1693;
    input [15:0] input_1694;
    input [15:0] input_1695;
    input [15:0] input_1696;
    input [15:0] input_1697;
    input [15:0] input_1698;
    input [15:0] input_1699;
    input [15:0] input_1700;
    input [15:0] input_1701;
    input [15:0] input_1702;
    input [15:0] input_1703;
    input [15:0] input_1704;
    input [15:0] input_1705;
    input [15:0] input_1706;
    input [15:0] input_1707;
    input [15:0] input_1708;
    input [15:0] input_1709;
    input [15:0] input_1710;
    input [15:0] input_1711;
    input [15:0] input_1712;
    input [15:0] input_1713;
    input [15:0] input_1714;
    input [15:0] input_1715;
    input [15:0] input_1716;
    input [15:0] input_1717;
    input [15:0] input_1718;
    input [15:0] input_1719;
    input [15:0] input_1720;
    input [15:0] input_1721;
    input [15:0] input_1722;
    input [15:0] input_1723;
    input [15:0] input_1724;
    input [15:0] input_1725;
    input [15:0] input_1726;
    input [15:0] input_1727;
    input [15:0] input_1728;
    input [15:0] input_1729;
    input [15:0] input_1730;
    input [15:0] input_1731;
    input [15:0] input_1732;
    input [15:0] input_1733;
    input [15:0] input_1734;
    input [15:0] input_1735;
    input [15:0] input_1736;
    input [15:0] input_1737;
    input [15:0] input_1738;
    input [15:0] input_1739;
    input [15:0] input_1740;
    input [15:0] input_1741;
    input [15:0] input_1742;
    input [15:0] input_1743;
    input [15:0] input_1744;
    input [15:0] input_1745;
    input [15:0] input_1746;
    input [15:0] input_1747;
    input [15:0] input_1748;
    input [15:0] input_1749;
    input [15:0] input_1750;
    input [15:0] input_1751;
    input [15:0] input_1752;
    input [15:0] input_1753;
    input [15:0] input_1754;
    input [15:0] input_1755;
    input [15:0] input_1756;
    input [15:0] input_1757;
    input [15:0] input_1758;
    input [15:0] input_1759;
    input [15:0] input_1760;
    input [15:0] input_1761;
    input [15:0] input_1762;
    input [15:0] input_1763;
    input [15:0] input_1764;
    input [15:0] input_1765;
    input [15:0] input_1766;
    input [15:0] input_1767;
    input [15:0] input_1768;
    input [15:0] input_1769;
    input [15:0] input_1770;
    input [15:0] input_1771;
    input [15:0] input_1772;
    input [15:0] input_1773;
    input [15:0] input_1774;
    input [15:0] input_1775;
    input [15:0] input_1776;
    input [15:0] input_1777;
    input [15:0] input_1778;
    input [15:0] input_1779;
    input [15:0] input_1780;
    input [15:0] input_1781;
    input [15:0] input_1782;
    input [15:0] input_1783;
    input [15:0] input_1784;
    input [15:0] input_1785;
    input [15:0] input_1786;
    input [15:0] input_1787;
    input [15:0] input_1788;
    input [15:0] input_1789;
    input [15:0] input_1790;
    input [15:0] input_1791;
    input [10:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      11'b00000000000 : begin
        result = input_0;
      end
      11'b00000000001 : begin
        result = input_1;
      end
      11'b00000000010 : begin
        result = input_2;
      end
      11'b00000000011 : begin
        result = input_3;
      end
      11'b00000000100 : begin
        result = input_4;
      end
      11'b00000000101 : begin
        result = input_5;
      end
      11'b00000000110 : begin
        result = input_6;
      end
      11'b00000000111 : begin
        result = input_7;
      end
      11'b00000001000 : begin
        result = input_8;
      end
      11'b00000001001 : begin
        result = input_9;
      end
      11'b00000001010 : begin
        result = input_10;
      end
      11'b00000001011 : begin
        result = input_11;
      end
      11'b00000001100 : begin
        result = input_12;
      end
      11'b00000001101 : begin
        result = input_13;
      end
      11'b00000001110 : begin
        result = input_14;
      end
      11'b00000001111 : begin
        result = input_15;
      end
      11'b00000010000 : begin
        result = input_16;
      end
      11'b00000010001 : begin
        result = input_17;
      end
      11'b00000010010 : begin
        result = input_18;
      end
      11'b00000010011 : begin
        result = input_19;
      end
      11'b00000010100 : begin
        result = input_20;
      end
      11'b00000010101 : begin
        result = input_21;
      end
      11'b00000010110 : begin
        result = input_22;
      end
      11'b00000010111 : begin
        result = input_23;
      end
      11'b00000011000 : begin
        result = input_24;
      end
      11'b00000011001 : begin
        result = input_25;
      end
      11'b00000011010 : begin
        result = input_26;
      end
      11'b00000011011 : begin
        result = input_27;
      end
      11'b00000011100 : begin
        result = input_28;
      end
      11'b00000011101 : begin
        result = input_29;
      end
      11'b00000011110 : begin
        result = input_30;
      end
      11'b00000011111 : begin
        result = input_31;
      end
      11'b00000100000 : begin
        result = input_32;
      end
      11'b00000100001 : begin
        result = input_33;
      end
      11'b00000100010 : begin
        result = input_34;
      end
      11'b00000100011 : begin
        result = input_35;
      end
      11'b00000100100 : begin
        result = input_36;
      end
      11'b00000100101 : begin
        result = input_37;
      end
      11'b00000100110 : begin
        result = input_38;
      end
      11'b00000100111 : begin
        result = input_39;
      end
      11'b00000101000 : begin
        result = input_40;
      end
      11'b00000101001 : begin
        result = input_41;
      end
      11'b00000101010 : begin
        result = input_42;
      end
      11'b00000101011 : begin
        result = input_43;
      end
      11'b00000101100 : begin
        result = input_44;
      end
      11'b00000101101 : begin
        result = input_45;
      end
      11'b00000101110 : begin
        result = input_46;
      end
      11'b00000101111 : begin
        result = input_47;
      end
      11'b00000110000 : begin
        result = input_48;
      end
      11'b00000110001 : begin
        result = input_49;
      end
      11'b00000110010 : begin
        result = input_50;
      end
      11'b00000110011 : begin
        result = input_51;
      end
      11'b00000110100 : begin
        result = input_52;
      end
      11'b00000110101 : begin
        result = input_53;
      end
      11'b00000110110 : begin
        result = input_54;
      end
      11'b00000110111 : begin
        result = input_55;
      end
      11'b00000111000 : begin
        result = input_56;
      end
      11'b00000111001 : begin
        result = input_57;
      end
      11'b00000111010 : begin
        result = input_58;
      end
      11'b00000111011 : begin
        result = input_59;
      end
      11'b00000111100 : begin
        result = input_60;
      end
      11'b00000111101 : begin
        result = input_61;
      end
      11'b00000111110 : begin
        result = input_62;
      end
      11'b00000111111 : begin
        result = input_63;
      end
      11'b00001000000 : begin
        result = input_64;
      end
      11'b00001000001 : begin
        result = input_65;
      end
      11'b00001000010 : begin
        result = input_66;
      end
      11'b00001000011 : begin
        result = input_67;
      end
      11'b00001000100 : begin
        result = input_68;
      end
      11'b00001000101 : begin
        result = input_69;
      end
      11'b00001000110 : begin
        result = input_70;
      end
      11'b00001000111 : begin
        result = input_71;
      end
      11'b00001001000 : begin
        result = input_72;
      end
      11'b00001001001 : begin
        result = input_73;
      end
      11'b00001001010 : begin
        result = input_74;
      end
      11'b00001001011 : begin
        result = input_75;
      end
      11'b00001001100 : begin
        result = input_76;
      end
      11'b00001001101 : begin
        result = input_77;
      end
      11'b00001001110 : begin
        result = input_78;
      end
      11'b00001001111 : begin
        result = input_79;
      end
      11'b00001010000 : begin
        result = input_80;
      end
      11'b00001010001 : begin
        result = input_81;
      end
      11'b00001010010 : begin
        result = input_82;
      end
      11'b00001010011 : begin
        result = input_83;
      end
      11'b00001010100 : begin
        result = input_84;
      end
      11'b00001010101 : begin
        result = input_85;
      end
      11'b00001010110 : begin
        result = input_86;
      end
      11'b00001010111 : begin
        result = input_87;
      end
      11'b00001011000 : begin
        result = input_88;
      end
      11'b00001011001 : begin
        result = input_89;
      end
      11'b00001011010 : begin
        result = input_90;
      end
      11'b00001011011 : begin
        result = input_91;
      end
      11'b00001011100 : begin
        result = input_92;
      end
      11'b00001011101 : begin
        result = input_93;
      end
      11'b00001011110 : begin
        result = input_94;
      end
      11'b00001011111 : begin
        result = input_95;
      end
      11'b00001100000 : begin
        result = input_96;
      end
      11'b00001100001 : begin
        result = input_97;
      end
      11'b00001100010 : begin
        result = input_98;
      end
      11'b00001100011 : begin
        result = input_99;
      end
      11'b00001100100 : begin
        result = input_100;
      end
      11'b00001100101 : begin
        result = input_101;
      end
      11'b00001100110 : begin
        result = input_102;
      end
      11'b00001100111 : begin
        result = input_103;
      end
      11'b00001101000 : begin
        result = input_104;
      end
      11'b00001101001 : begin
        result = input_105;
      end
      11'b00001101010 : begin
        result = input_106;
      end
      11'b00001101011 : begin
        result = input_107;
      end
      11'b00001101100 : begin
        result = input_108;
      end
      11'b00001101101 : begin
        result = input_109;
      end
      11'b00001101110 : begin
        result = input_110;
      end
      11'b00001101111 : begin
        result = input_111;
      end
      11'b00001110000 : begin
        result = input_112;
      end
      11'b00001110001 : begin
        result = input_113;
      end
      11'b00001110010 : begin
        result = input_114;
      end
      11'b00001110011 : begin
        result = input_115;
      end
      11'b00001110100 : begin
        result = input_116;
      end
      11'b00001110101 : begin
        result = input_117;
      end
      11'b00001110110 : begin
        result = input_118;
      end
      11'b00001110111 : begin
        result = input_119;
      end
      11'b00001111000 : begin
        result = input_120;
      end
      11'b00001111001 : begin
        result = input_121;
      end
      11'b00001111010 : begin
        result = input_122;
      end
      11'b00001111011 : begin
        result = input_123;
      end
      11'b00001111100 : begin
        result = input_124;
      end
      11'b00001111101 : begin
        result = input_125;
      end
      11'b00001111110 : begin
        result = input_126;
      end
      11'b00001111111 : begin
        result = input_127;
      end
      11'b00010000000 : begin
        result = input_128;
      end
      11'b00010000001 : begin
        result = input_129;
      end
      11'b00010000010 : begin
        result = input_130;
      end
      11'b00010000011 : begin
        result = input_131;
      end
      11'b00010000100 : begin
        result = input_132;
      end
      11'b00010000101 : begin
        result = input_133;
      end
      11'b00010000110 : begin
        result = input_134;
      end
      11'b00010000111 : begin
        result = input_135;
      end
      11'b00010001000 : begin
        result = input_136;
      end
      11'b00010001001 : begin
        result = input_137;
      end
      11'b00010001010 : begin
        result = input_138;
      end
      11'b00010001011 : begin
        result = input_139;
      end
      11'b00010001100 : begin
        result = input_140;
      end
      11'b00010001101 : begin
        result = input_141;
      end
      11'b00010001110 : begin
        result = input_142;
      end
      11'b00010001111 : begin
        result = input_143;
      end
      11'b00010010000 : begin
        result = input_144;
      end
      11'b00010010001 : begin
        result = input_145;
      end
      11'b00010010010 : begin
        result = input_146;
      end
      11'b00010010011 : begin
        result = input_147;
      end
      11'b00010010100 : begin
        result = input_148;
      end
      11'b00010010101 : begin
        result = input_149;
      end
      11'b00010010110 : begin
        result = input_150;
      end
      11'b00010010111 : begin
        result = input_151;
      end
      11'b00010011000 : begin
        result = input_152;
      end
      11'b00010011001 : begin
        result = input_153;
      end
      11'b00010011010 : begin
        result = input_154;
      end
      11'b00010011011 : begin
        result = input_155;
      end
      11'b00010011100 : begin
        result = input_156;
      end
      11'b00010011101 : begin
        result = input_157;
      end
      11'b00010011110 : begin
        result = input_158;
      end
      11'b00010011111 : begin
        result = input_159;
      end
      11'b00010100000 : begin
        result = input_160;
      end
      11'b00010100001 : begin
        result = input_161;
      end
      11'b00010100010 : begin
        result = input_162;
      end
      11'b00010100011 : begin
        result = input_163;
      end
      11'b00010100100 : begin
        result = input_164;
      end
      11'b00010100101 : begin
        result = input_165;
      end
      11'b00010100110 : begin
        result = input_166;
      end
      11'b00010100111 : begin
        result = input_167;
      end
      11'b00010101000 : begin
        result = input_168;
      end
      11'b00010101001 : begin
        result = input_169;
      end
      11'b00010101010 : begin
        result = input_170;
      end
      11'b00010101011 : begin
        result = input_171;
      end
      11'b00010101100 : begin
        result = input_172;
      end
      11'b00010101101 : begin
        result = input_173;
      end
      11'b00010101110 : begin
        result = input_174;
      end
      11'b00010101111 : begin
        result = input_175;
      end
      11'b00010110000 : begin
        result = input_176;
      end
      11'b00010110001 : begin
        result = input_177;
      end
      11'b00010110010 : begin
        result = input_178;
      end
      11'b00010110011 : begin
        result = input_179;
      end
      11'b00010110100 : begin
        result = input_180;
      end
      11'b00010110101 : begin
        result = input_181;
      end
      11'b00010110110 : begin
        result = input_182;
      end
      11'b00010110111 : begin
        result = input_183;
      end
      11'b00010111000 : begin
        result = input_184;
      end
      11'b00010111001 : begin
        result = input_185;
      end
      11'b00010111010 : begin
        result = input_186;
      end
      11'b00010111011 : begin
        result = input_187;
      end
      11'b00010111100 : begin
        result = input_188;
      end
      11'b00010111101 : begin
        result = input_189;
      end
      11'b00010111110 : begin
        result = input_190;
      end
      11'b00010111111 : begin
        result = input_191;
      end
      11'b00011000000 : begin
        result = input_192;
      end
      11'b00011000001 : begin
        result = input_193;
      end
      11'b00011000010 : begin
        result = input_194;
      end
      11'b00011000011 : begin
        result = input_195;
      end
      11'b00011000100 : begin
        result = input_196;
      end
      11'b00011000101 : begin
        result = input_197;
      end
      11'b00011000110 : begin
        result = input_198;
      end
      11'b00011000111 : begin
        result = input_199;
      end
      11'b00011001000 : begin
        result = input_200;
      end
      11'b00011001001 : begin
        result = input_201;
      end
      11'b00011001010 : begin
        result = input_202;
      end
      11'b00011001011 : begin
        result = input_203;
      end
      11'b00011001100 : begin
        result = input_204;
      end
      11'b00011001101 : begin
        result = input_205;
      end
      11'b00011001110 : begin
        result = input_206;
      end
      11'b00011001111 : begin
        result = input_207;
      end
      11'b00011010000 : begin
        result = input_208;
      end
      11'b00011010001 : begin
        result = input_209;
      end
      11'b00011010010 : begin
        result = input_210;
      end
      11'b00011010011 : begin
        result = input_211;
      end
      11'b00011010100 : begin
        result = input_212;
      end
      11'b00011010101 : begin
        result = input_213;
      end
      11'b00011010110 : begin
        result = input_214;
      end
      11'b00011010111 : begin
        result = input_215;
      end
      11'b00011011000 : begin
        result = input_216;
      end
      11'b00011011001 : begin
        result = input_217;
      end
      11'b00011011010 : begin
        result = input_218;
      end
      11'b00011011011 : begin
        result = input_219;
      end
      11'b00011011100 : begin
        result = input_220;
      end
      11'b00011011101 : begin
        result = input_221;
      end
      11'b00011011110 : begin
        result = input_222;
      end
      11'b00011011111 : begin
        result = input_223;
      end
      11'b00011100000 : begin
        result = input_224;
      end
      11'b00011100001 : begin
        result = input_225;
      end
      11'b00011100010 : begin
        result = input_226;
      end
      11'b00011100011 : begin
        result = input_227;
      end
      11'b00011100100 : begin
        result = input_228;
      end
      11'b00011100101 : begin
        result = input_229;
      end
      11'b00011100110 : begin
        result = input_230;
      end
      11'b00011100111 : begin
        result = input_231;
      end
      11'b00011101000 : begin
        result = input_232;
      end
      11'b00011101001 : begin
        result = input_233;
      end
      11'b00011101010 : begin
        result = input_234;
      end
      11'b00011101011 : begin
        result = input_235;
      end
      11'b00011101100 : begin
        result = input_236;
      end
      11'b00011101101 : begin
        result = input_237;
      end
      11'b00011101110 : begin
        result = input_238;
      end
      11'b00011101111 : begin
        result = input_239;
      end
      11'b00011110000 : begin
        result = input_240;
      end
      11'b00011110001 : begin
        result = input_241;
      end
      11'b00011110010 : begin
        result = input_242;
      end
      11'b00011110011 : begin
        result = input_243;
      end
      11'b00011110100 : begin
        result = input_244;
      end
      11'b00011110101 : begin
        result = input_245;
      end
      11'b00011110110 : begin
        result = input_246;
      end
      11'b00011110111 : begin
        result = input_247;
      end
      11'b00011111000 : begin
        result = input_248;
      end
      11'b00011111001 : begin
        result = input_249;
      end
      11'b00011111010 : begin
        result = input_250;
      end
      11'b00011111011 : begin
        result = input_251;
      end
      11'b00011111100 : begin
        result = input_252;
      end
      11'b00011111101 : begin
        result = input_253;
      end
      11'b00011111110 : begin
        result = input_254;
      end
      11'b00011111111 : begin
        result = input_255;
      end
      11'b00100000000 : begin
        result = input_256;
      end
      11'b00100000001 : begin
        result = input_257;
      end
      11'b00100000010 : begin
        result = input_258;
      end
      11'b00100000011 : begin
        result = input_259;
      end
      11'b00100000100 : begin
        result = input_260;
      end
      11'b00100000101 : begin
        result = input_261;
      end
      11'b00100000110 : begin
        result = input_262;
      end
      11'b00100000111 : begin
        result = input_263;
      end
      11'b00100001000 : begin
        result = input_264;
      end
      11'b00100001001 : begin
        result = input_265;
      end
      11'b00100001010 : begin
        result = input_266;
      end
      11'b00100001011 : begin
        result = input_267;
      end
      11'b00100001100 : begin
        result = input_268;
      end
      11'b00100001101 : begin
        result = input_269;
      end
      11'b00100001110 : begin
        result = input_270;
      end
      11'b00100001111 : begin
        result = input_271;
      end
      11'b00100010000 : begin
        result = input_272;
      end
      11'b00100010001 : begin
        result = input_273;
      end
      11'b00100010010 : begin
        result = input_274;
      end
      11'b00100010011 : begin
        result = input_275;
      end
      11'b00100010100 : begin
        result = input_276;
      end
      11'b00100010101 : begin
        result = input_277;
      end
      11'b00100010110 : begin
        result = input_278;
      end
      11'b00100010111 : begin
        result = input_279;
      end
      11'b00100011000 : begin
        result = input_280;
      end
      11'b00100011001 : begin
        result = input_281;
      end
      11'b00100011010 : begin
        result = input_282;
      end
      11'b00100011011 : begin
        result = input_283;
      end
      11'b00100011100 : begin
        result = input_284;
      end
      11'b00100011101 : begin
        result = input_285;
      end
      11'b00100011110 : begin
        result = input_286;
      end
      11'b00100011111 : begin
        result = input_287;
      end
      11'b00100100000 : begin
        result = input_288;
      end
      11'b00100100001 : begin
        result = input_289;
      end
      11'b00100100010 : begin
        result = input_290;
      end
      11'b00100100011 : begin
        result = input_291;
      end
      11'b00100100100 : begin
        result = input_292;
      end
      11'b00100100101 : begin
        result = input_293;
      end
      11'b00100100110 : begin
        result = input_294;
      end
      11'b00100100111 : begin
        result = input_295;
      end
      11'b00100101000 : begin
        result = input_296;
      end
      11'b00100101001 : begin
        result = input_297;
      end
      11'b00100101010 : begin
        result = input_298;
      end
      11'b00100101011 : begin
        result = input_299;
      end
      11'b00100101100 : begin
        result = input_300;
      end
      11'b00100101101 : begin
        result = input_301;
      end
      11'b00100101110 : begin
        result = input_302;
      end
      11'b00100101111 : begin
        result = input_303;
      end
      11'b00100110000 : begin
        result = input_304;
      end
      11'b00100110001 : begin
        result = input_305;
      end
      11'b00100110010 : begin
        result = input_306;
      end
      11'b00100110011 : begin
        result = input_307;
      end
      11'b00100110100 : begin
        result = input_308;
      end
      11'b00100110101 : begin
        result = input_309;
      end
      11'b00100110110 : begin
        result = input_310;
      end
      11'b00100110111 : begin
        result = input_311;
      end
      11'b00100111000 : begin
        result = input_312;
      end
      11'b00100111001 : begin
        result = input_313;
      end
      11'b00100111010 : begin
        result = input_314;
      end
      11'b00100111011 : begin
        result = input_315;
      end
      11'b00100111100 : begin
        result = input_316;
      end
      11'b00100111101 : begin
        result = input_317;
      end
      11'b00100111110 : begin
        result = input_318;
      end
      11'b00100111111 : begin
        result = input_319;
      end
      11'b00101000000 : begin
        result = input_320;
      end
      11'b00101000001 : begin
        result = input_321;
      end
      11'b00101000010 : begin
        result = input_322;
      end
      11'b00101000011 : begin
        result = input_323;
      end
      11'b00101000100 : begin
        result = input_324;
      end
      11'b00101000101 : begin
        result = input_325;
      end
      11'b00101000110 : begin
        result = input_326;
      end
      11'b00101000111 : begin
        result = input_327;
      end
      11'b00101001000 : begin
        result = input_328;
      end
      11'b00101001001 : begin
        result = input_329;
      end
      11'b00101001010 : begin
        result = input_330;
      end
      11'b00101001011 : begin
        result = input_331;
      end
      11'b00101001100 : begin
        result = input_332;
      end
      11'b00101001101 : begin
        result = input_333;
      end
      11'b00101001110 : begin
        result = input_334;
      end
      11'b00101001111 : begin
        result = input_335;
      end
      11'b00101010000 : begin
        result = input_336;
      end
      11'b00101010001 : begin
        result = input_337;
      end
      11'b00101010010 : begin
        result = input_338;
      end
      11'b00101010011 : begin
        result = input_339;
      end
      11'b00101010100 : begin
        result = input_340;
      end
      11'b00101010101 : begin
        result = input_341;
      end
      11'b00101010110 : begin
        result = input_342;
      end
      11'b00101010111 : begin
        result = input_343;
      end
      11'b00101011000 : begin
        result = input_344;
      end
      11'b00101011001 : begin
        result = input_345;
      end
      11'b00101011010 : begin
        result = input_346;
      end
      11'b00101011011 : begin
        result = input_347;
      end
      11'b00101011100 : begin
        result = input_348;
      end
      11'b00101011101 : begin
        result = input_349;
      end
      11'b00101011110 : begin
        result = input_350;
      end
      11'b00101011111 : begin
        result = input_351;
      end
      11'b00101100000 : begin
        result = input_352;
      end
      11'b00101100001 : begin
        result = input_353;
      end
      11'b00101100010 : begin
        result = input_354;
      end
      11'b00101100011 : begin
        result = input_355;
      end
      11'b00101100100 : begin
        result = input_356;
      end
      11'b00101100101 : begin
        result = input_357;
      end
      11'b00101100110 : begin
        result = input_358;
      end
      11'b00101100111 : begin
        result = input_359;
      end
      11'b00101101000 : begin
        result = input_360;
      end
      11'b00101101001 : begin
        result = input_361;
      end
      11'b00101101010 : begin
        result = input_362;
      end
      11'b00101101011 : begin
        result = input_363;
      end
      11'b00101101100 : begin
        result = input_364;
      end
      11'b00101101101 : begin
        result = input_365;
      end
      11'b00101101110 : begin
        result = input_366;
      end
      11'b00101101111 : begin
        result = input_367;
      end
      11'b00101110000 : begin
        result = input_368;
      end
      11'b00101110001 : begin
        result = input_369;
      end
      11'b00101110010 : begin
        result = input_370;
      end
      11'b00101110011 : begin
        result = input_371;
      end
      11'b00101110100 : begin
        result = input_372;
      end
      11'b00101110101 : begin
        result = input_373;
      end
      11'b00101110110 : begin
        result = input_374;
      end
      11'b00101110111 : begin
        result = input_375;
      end
      11'b00101111000 : begin
        result = input_376;
      end
      11'b00101111001 : begin
        result = input_377;
      end
      11'b00101111010 : begin
        result = input_378;
      end
      11'b00101111011 : begin
        result = input_379;
      end
      11'b00101111100 : begin
        result = input_380;
      end
      11'b00101111101 : begin
        result = input_381;
      end
      11'b00101111110 : begin
        result = input_382;
      end
      11'b00101111111 : begin
        result = input_383;
      end
      11'b00110000000 : begin
        result = input_384;
      end
      11'b00110000001 : begin
        result = input_385;
      end
      11'b00110000010 : begin
        result = input_386;
      end
      11'b00110000011 : begin
        result = input_387;
      end
      11'b00110000100 : begin
        result = input_388;
      end
      11'b00110000101 : begin
        result = input_389;
      end
      11'b00110000110 : begin
        result = input_390;
      end
      11'b00110000111 : begin
        result = input_391;
      end
      11'b00110001000 : begin
        result = input_392;
      end
      11'b00110001001 : begin
        result = input_393;
      end
      11'b00110001010 : begin
        result = input_394;
      end
      11'b00110001011 : begin
        result = input_395;
      end
      11'b00110001100 : begin
        result = input_396;
      end
      11'b00110001101 : begin
        result = input_397;
      end
      11'b00110001110 : begin
        result = input_398;
      end
      11'b00110001111 : begin
        result = input_399;
      end
      11'b00110010000 : begin
        result = input_400;
      end
      11'b00110010001 : begin
        result = input_401;
      end
      11'b00110010010 : begin
        result = input_402;
      end
      11'b00110010011 : begin
        result = input_403;
      end
      11'b00110010100 : begin
        result = input_404;
      end
      11'b00110010101 : begin
        result = input_405;
      end
      11'b00110010110 : begin
        result = input_406;
      end
      11'b00110010111 : begin
        result = input_407;
      end
      11'b00110011000 : begin
        result = input_408;
      end
      11'b00110011001 : begin
        result = input_409;
      end
      11'b00110011010 : begin
        result = input_410;
      end
      11'b00110011011 : begin
        result = input_411;
      end
      11'b00110011100 : begin
        result = input_412;
      end
      11'b00110011101 : begin
        result = input_413;
      end
      11'b00110011110 : begin
        result = input_414;
      end
      11'b00110011111 : begin
        result = input_415;
      end
      11'b00110100000 : begin
        result = input_416;
      end
      11'b00110100001 : begin
        result = input_417;
      end
      11'b00110100010 : begin
        result = input_418;
      end
      11'b00110100011 : begin
        result = input_419;
      end
      11'b00110100100 : begin
        result = input_420;
      end
      11'b00110100101 : begin
        result = input_421;
      end
      11'b00110100110 : begin
        result = input_422;
      end
      11'b00110100111 : begin
        result = input_423;
      end
      11'b00110101000 : begin
        result = input_424;
      end
      11'b00110101001 : begin
        result = input_425;
      end
      11'b00110101010 : begin
        result = input_426;
      end
      11'b00110101011 : begin
        result = input_427;
      end
      11'b00110101100 : begin
        result = input_428;
      end
      11'b00110101101 : begin
        result = input_429;
      end
      11'b00110101110 : begin
        result = input_430;
      end
      11'b00110101111 : begin
        result = input_431;
      end
      11'b00110110000 : begin
        result = input_432;
      end
      11'b00110110001 : begin
        result = input_433;
      end
      11'b00110110010 : begin
        result = input_434;
      end
      11'b00110110011 : begin
        result = input_435;
      end
      11'b00110110100 : begin
        result = input_436;
      end
      11'b00110110101 : begin
        result = input_437;
      end
      11'b00110110110 : begin
        result = input_438;
      end
      11'b00110110111 : begin
        result = input_439;
      end
      11'b00110111000 : begin
        result = input_440;
      end
      11'b00110111001 : begin
        result = input_441;
      end
      11'b00110111010 : begin
        result = input_442;
      end
      11'b00110111011 : begin
        result = input_443;
      end
      11'b00110111100 : begin
        result = input_444;
      end
      11'b00110111101 : begin
        result = input_445;
      end
      11'b00110111110 : begin
        result = input_446;
      end
      11'b00110111111 : begin
        result = input_447;
      end
      11'b00111000000 : begin
        result = input_448;
      end
      11'b00111000001 : begin
        result = input_449;
      end
      11'b00111000010 : begin
        result = input_450;
      end
      11'b00111000011 : begin
        result = input_451;
      end
      11'b00111000100 : begin
        result = input_452;
      end
      11'b00111000101 : begin
        result = input_453;
      end
      11'b00111000110 : begin
        result = input_454;
      end
      11'b00111000111 : begin
        result = input_455;
      end
      11'b00111001000 : begin
        result = input_456;
      end
      11'b00111001001 : begin
        result = input_457;
      end
      11'b00111001010 : begin
        result = input_458;
      end
      11'b00111001011 : begin
        result = input_459;
      end
      11'b00111001100 : begin
        result = input_460;
      end
      11'b00111001101 : begin
        result = input_461;
      end
      11'b00111001110 : begin
        result = input_462;
      end
      11'b00111001111 : begin
        result = input_463;
      end
      11'b00111010000 : begin
        result = input_464;
      end
      11'b00111010001 : begin
        result = input_465;
      end
      11'b00111010010 : begin
        result = input_466;
      end
      11'b00111010011 : begin
        result = input_467;
      end
      11'b00111010100 : begin
        result = input_468;
      end
      11'b00111010101 : begin
        result = input_469;
      end
      11'b00111010110 : begin
        result = input_470;
      end
      11'b00111010111 : begin
        result = input_471;
      end
      11'b00111011000 : begin
        result = input_472;
      end
      11'b00111011001 : begin
        result = input_473;
      end
      11'b00111011010 : begin
        result = input_474;
      end
      11'b00111011011 : begin
        result = input_475;
      end
      11'b00111011100 : begin
        result = input_476;
      end
      11'b00111011101 : begin
        result = input_477;
      end
      11'b00111011110 : begin
        result = input_478;
      end
      11'b00111011111 : begin
        result = input_479;
      end
      11'b00111100000 : begin
        result = input_480;
      end
      11'b00111100001 : begin
        result = input_481;
      end
      11'b00111100010 : begin
        result = input_482;
      end
      11'b00111100011 : begin
        result = input_483;
      end
      11'b00111100100 : begin
        result = input_484;
      end
      11'b00111100101 : begin
        result = input_485;
      end
      11'b00111100110 : begin
        result = input_486;
      end
      11'b00111100111 : begin
        result = input_487;
      end
      11'b00111101000 : begin
        result = input_488;
      end
      11'b00111101001 : begin
        result = input_489;
      end
      11'b00111101010 : begin
        result = input_490;
      end
      11'b00111101011 : begin
        result = input_491;
      end
      11'b00111101100 : begin
        result = input_492;
      end
      11'b00111101101 : begin
        result = input_493;
      end
      11'b00111101110 : begin
        result = input_494;
      end
      11'b00111101111 : begin
        result = input_495;
      end
      11'b00111110000 : begin
        result = input_496;
      end
      11'b00111110001 : begin
        result = input_497;
      end
      11'b00111110010 : begin
        result = input_498;
      end
      11'b00111110011 : begin
        result = input_499;
      end
      11'b00111110100 : begin
        result = input_500;
      end
      11'b00111110101 : begin
        result = input_501;
      end
      11'b00111110110 : begin
        result = input_502;
      end
      11'b00111110111 : begin
        result = input_503;
      end
      11'b00111111000 : begin
        result = input_504;
      end
      11'b00111111001 : begin
        result = input_505;
      end
      11'b00111111010 : begin
        result = input_506;
      end
      11'b00111111011 : begin
        result = input_507;
      end
      11'b00111111100 : begin
        result = input_508;
      end
      11'b00111111101 : begin
        result = input_509;
      end
      11'b00111111110 : begin
        result = input_510;
      end
      11'b00111111111 : begin
        result = input_511;
      end
      11'b01000000000 : begin
        result = input_512;
      end
      11'b01000000001 : begin
        result = input_513;
      end
      11'b01000000010 : begin
        result = input_514;
      end
      11'b01000000011 : begin
        result = input_515;
      end
      11'b01000000100 : begin
        result = input_516;
      end
      11'b01000000101 : begin
        result = input_517;
      end
      11'b01000000110 : begin
        result = input_518;
      end
      11'b01000000111 : begin
        result = input_519;
      end
      11'b01000001000 : begin
        result = input_520;
      end
      11'b01000001001 : begin
        result = input_521;
      end
      11'b01000001010 : begin
        result = input_522;
      end
      11'b01000001011 : begin
        result = input_523;
      end
      11'b01000001100 : begin
        result = input_524;
      end
      11'b01000001101 : begin
        result = input_525;
      end
      11'b01000001110 : begin
        result = input_526;
      end
      11'b01000001111 : begin
        result = input_527;
      end
      11'b01000010000 : begin
        result = input_528;
      end
      11'b01000010001 : begin
        result = input_529;
      end
      11'b01000010010 : begin
        result = input_530;
      end
      11'b01000010011 : begin
        result = input_531;
      end
      11'b01000010100 : begin
        result = input_532;
      end
      11'b01000010101 : begin
        result = input_533;
      end
      11'b01000010110 : begin
        result = input_534;
      end
      11'b01000010111 : begin
        result = input_535;
      end
      11'b01000011000 : begin
        result = input_536;
      end
      11'b01000011001 : begin
        result = input_537;
      end
      11'b01000011010 : begin
        result = input_538;
      end
      11'b01000011011 : begin
        result = input_539;
      end
      11'b01000011100 : begin
        result = input_540;
      end
      11'b01000011101 : begin
        result = input_541;
      end
      11'b01000011110 : begin
        result = input_542;
      end
      11'b01000011111 : begin
        result = input_543;
      end
      11'b01000100000 : begin
        result = input_544;
      end
      11'b01000100001 : begin
        result = input_545;
      end
      11'b01000100010 : begin
        result = input_546;
      end
      11'b01000100011 : begin
        result = input_547;
      end
      11'b01000100100 : begin
        result = input_548;
      end
      11'b01000100101 : begin
        result = input_549;
      end
      11'b01000100110 : begin
        result = input_550;
      end
      11'b01000100111 : begin
        result = input_551;
      end
      11'b01000101000 : begin
        result = input_552;
      end
      11'b01000101001 : begin
        result = input_553;
      end
      11'b01000101010 : begin
        result = input_554;
      end
      11'b01000101011 : begin
        result = input_555;
      end
      11'b01000101100 : begin
        result = input_556;
      end
      11'b01000101101 : begin
        result = input_557;
      end
      11'b01000101110 : begin
        result = input_558;
      end
      11'b01000101111 : begin
        result = input_559;
      end
      11'b01000110000 : begin
        result = input_560;
      end
      11'b01000110001 : begin
        result = input_561;
      end
      11'b01000110010 : begin
        result = input_562;
      end
      11'b01000110011 : begin
        result = input_563;
      end
      11'b01000110100 : begin
        result = input_564;
      end
      11'b01000110101 : begin
        result = input_565;
      end
      11'b01000110110 : begin
        result = input_566;
      end
      11'b01000110111 : begin
        result = input_567;
      end
      11'b01000111000 : begin
        result = input_568;
      end
      11'b01000111001 : begin
        result = input_569;
      end
      11'b01000111010 : begin
        result = input_570;
      end
      11'b01000111011 : begin
        result = input_571;
      end
      11'b01000111100 : begin
        result = input_572;
      end
      11'b01000111101 : begin
        result = input_573;
      end
      11'b01000111110 : begin
        result = input_574;
      end
      11'b01000111111 : begin
        result = input_575;
      end
      11'b01001000000 : begin
        result = input_576;
      end
      11'b01001000001 : begin
        result = input_577;
      end
      11'b01001000010 : begin
        result = input_578;
      end
      11'b01001000011 : begin
        result = input_579;
      end
      11'b01001000100 : begin
        result = input_580;
      end
      11'b01001000101 : begin
        result = input_581;
      end
      11'b01001000110 : begin
        result = input_582;
      end
      11'b01001000111 : begin
        result = input_583;
      end
      11'b01001001000 : begin
        result = input_584;
      end
      11'b01001001001 : begin
        result = input_585;
      end
      11'b01001001010 : begin
        result = input_586;
      end
      11'b01001001011 : begin
        result = input_587;
      end
      11'b01001001100 : begin
        result = input_588;
      end
      11'b01001001101 : begin
        result = input_589;
      end
      11'b01001001110 : begin
        result = input_590;
      end
      11'b01001001111 : begin
        result = input_591;
      end
      11'b01001010000 : begin
        result = input_592;
      end
      11'b01001010001 : begin
        result = input_593;
      end
      11'b01001010010 : begin
        result = input_594;
      end
      11'b01001010011 : begin
        result = input_595;
      end
      11'b01001010100 : begin
        result = input_596;
      end
      11'b01001010101 : begin
        result = input_597;
      end
      11'b01001010110 : begin
        result = input_598;
      end
      11'b01001010111 : begin
        result = input_599;
      end
      11'b01001011000 : begin
        result = input_600;
      end
      11'b01001011001 : begin
        result = input_601;
      end
      11'b01001011010 : begin
        result = input_602;
      end
      11'b01001011011 : begin
        result = input_603;
      end
      11'b01001011100 : begin
        result = input_604;
      end
      11'b01001011101 : begin
        result = input_605;
      end
      11'b01001011110 : begin
        result = input_606;
      end
      11'b01001011111 : begin
        result = input_607;
      end
      11'b01001100000 : begin
        result = input_608;
      end
      11'b01001100001 : begin
        result = input_609;
      end
      11'b01001100010 : begin
        result = input_610;
      end
      11'b01001100011 : begin
        result = input_611;
      end
      11'b01001100100 : begin
        result = input_612;
      end
      11'b01001100101 : begin
        result = input_613;
      end
      11'b01001100110 : begin
        result = input_614;
      end
      11'b01001100111 : begin
        result = input_615;
      end
      11'b01001101000 : begin
        result = input_616;
      end
      11'b01001101001 : begin
        result = input_617;
      end
      11'b01001101010 : begin
        result = input_618;
      end
      11'b01001101011 : begin
        result = input_619;
      end
      11'b01001101100 : begin
        result = input_620;
      end
      11'b01001101101 : begin
        result = input_621;
      end
      11'b01001101110 : begin
        result = input_622;
      end
      11'b01001101111 : begin
        result = input_623;
      end
      11'b01001110000 : begin
        result = input_624;
      end
      11'b01001110001 : begin
        result = input_625;
      end
      11'b01001110010 : begin
        result = input_626;
      end
      11'b01001110011 : begin
        result = input_627;
      end
      11'b01001110100 : begin
        result = input_628;
      end
      11'b01001110101 : begin
        result = input_629;
      end
      11'b01001110110 : begin
        result = input_630;
      end
      11'b01001110111 : begin
        result = input_631;
      end
      11'b01001111000 : begin
        result = input_632;
      end
      11'b01001111001 : begin
        result = input_633;
      end
      11'b01001111010 : begin
        result = input_634;
      end
      11'b01001111011 : begin
        result = input_635;
      end
      11'b01001111100 : begin
        result = input_636;
      end
      11'b01001111101 : begin
        result = input_637;
      end
      11'b01001111110 : begin
        result = input_638;
      end
      11'b01001111111 : begin
        result = input_639;
      end
      11'b01010000000 : begin
        result = input_640;
      end
      11'b01010000001 : begin
        result = input_641;
      end
      11'b01010000010 : begin
        result = input_642;
      end
      11'b01010000011 : begin
        result = input_643;
      end
      11'b01010000100 : begin
        result = input_644;
      end
      11'b01010000101 : begin
        result = input_645;
      end
      11'b01010000110 : begin
        result = input_646;
      end
      11'b01010000111 : begin
        result = input_647;
      end
      11'b01010001000 : begin
        result = input_648;
      end
      11'b01010001001 : begin
        result = input_649;
      end
      11'b01010001010 : begin
        result = input_650;
      end
      11'b01010001011 : begin
        result = input_651;
      end
      11'b01010001100 : begin
        result = input_652;
      end
      11'b01010001101 : begin
        result = input_653;
      end
      11'b01010001110 : begin
        result = input_654;
      end
      11'b01010001111 : begin
        result = input_655;
      end
      11'b01010010000 : begin
        result = input_656;
      end
      11'b01010010001 : begin
        result = input_657;
      end
      11'b01010010010 : begin
        result = input_658;
      end
      11'b01010010011 : begin
        result = input_659;
      end
      11'b01010010100 : begin
        result = input_660;
      end
      11'b01010010101 : begin
        result = input_661;
      end
      11'b01010010110 : begin
        result = input_662;
      end
      11'b01010010111 : begin
        result = input_663;
      end
      11'b01010011000 : begin
        result = input_664;
      end
      11'b01010011001 : begin
        result = input_665;
      end
      11'b01010011010 : begin
        result = input_666;
      end
      11'b01010011011 : begin
        result = input_667;
      end
      11'b01010011100 : begin
        result = input_668;
      end
      11'b01010011101 : begin
        result = input_669;
      end
      11'b01010011110 : begin
        result = input_670;
      end
      11'b01010011111 : begin
        result = input_671;
      end
      11'b01010100000 : begin
        result = input_672;
      end
      11'b01010100001 : begin
        result = input_673;
      end
      11'b01010100010 : begin
        result = input_674;
      end
      11'b01010100011 : begin
        result = input_675;
      end
      11'b01010100100 : begin
        result = input_676;
      end
      11'b01010100101 : begin
        result = input_677;
      end
      11'b01010100110 : begin
        result = input_678;
      end
      11'b01010100111 : begin
        result = input_679;
      end
      11'b01010101000 : begin
        result = input_680;
      end
      11'b01010101001 : begin
        result = input_681;
      end
      11'b01010101010 : begin
        result = input_682;
      end
      11'b01010101011 : begin
        result = input_683;
      end
      11'b01010101100 : begin
        result = input_684;
      end
      11'b01010101101 : begin
        result = input_685;
      end
      11'b01010101110 : begin
        result = input_686;
      end
      11'b01010101111 : begin
        result = input_687;
      end
      11'b01010110000 : begin
        result = input_688;
      end
      11'b01010110001 : begin
        result = input_689;
      end
      11'b01010110010 : begin
        result = input_690;
      end
      11'b01010110011 : begin
        result = input_691;
      end
      11'b01010110100 : begin
        result = input_692;
      end
      11'b01010110101 : begin
        result = input_693;
      end
      11'b01010110110 : begin
        result = input_694;
      end
      11'b01010110111 : begin
        result = input_695;
      end
      11'b01010111000 : begin
        result = input_696;
      end
      11'b01010111001 : begin
        result = input_697;
      end
      11'b01010111010 : begin
        result = input_698;
      end
      11'b01010111011 : begin
        result = input_699;
      end
      11'b01010111100 : begin
        result = input_700;
      end
      11'b01010111101 : begin
        result = input_701;
      end
      11'b01010111110 : begin
        result = input_702;
      end
      11'b01010111111 : begin
        result = input_703;
      end
      11'b01011000000 : begin
        result = input_704;
      end
      11'b01011000001 : begin
        result = input_705;
      end
      11'b01011000010 : begin
        result = input_706;
      end
      11'b01011000011 : begin
        result = input_707;
      end
      11'b01011000100 : begin
        result = input_708;
      end
      11'b01011000101 : begin
        result = input_709;
      end
      11'b01011000110 : begin
        result = input_710;
      end
      11'b01011000111 : begin
        result = input_711;
      end
      11'b01011001000 : begin
        result = input_712;
      end
      11'b01011001001 : begin
        result = input_713;
      end
      11'b01011001010 : begin
        result = input_714;
      end
      11'b01011001011 : begin
        result = input_715;
      end
      11'b01011001100 : begin
        result = input_716;
      end
      11'b01011001101 : begin
        result = input_717;
      end
      11'b01011001110 : begin
        result = input_718;
      end
      11'b01011001111 : begin
        result = input_719;
      end
      11'b01011010000 : begin
        result = input_720;
      end
      11'b01011010001 : begin
        result = input_721;
      end
      11'b01011010010 : begin
        result = input_722;
      end
      11'b01011010011 : begin
        result = input_723;
      end
      11'b01011010100 : begin
        result = input_724;
      end
      11'b01011010101 : begin
        result = input_725;
      end
      11'b01011010110 : begin
        result = input_726;
      end
      11'b01011010111 : begin
        result = input_727;
      end
      11'b01011011000 : begin
        result = input_728;
      end
      11'b01011011001 : begin
        result = input_729;
      end
      11'b01011011010 : begin
        result = input_730;
      end
      11'b01011011011 : begin
        result = input_731;
      end
      11'b01011011100 : begin
        result = input_732;
      end
      11'b01011011101 : begin
        result = input_733;
      end
      11'b01011011110 : begin
        result = input_734;
      end
      11'b01011011111 : begin
        result = input_735;
      end
      11'b01011100000 : begin
        result = input_736;
      end
      11'b01011100001 : begin
        result = input_737;
      end
      11'b01011100010 : begin
        result = input_738;
      end
      11'b01011100011 : begin
        result = input_739;
      end
      11'b01011100100 : begin
        result = input_740;
      end
      11'b01011100101 : begin
        result = input_741;
      end
      11'b01011100110 : begin
        result = input_742;
      end
      11'b01011100111 : begin
        result = input_743;
      end
      11'b01011101000 : begin
        result = input_744;
      end
      11'b01011101001 : begin
        result = input_745;
      end
      11'b01011101010 : begin
        result = input_746;
      end
      11'b01011101011 : begin
        result = input_747;
      end
      11'b01011101100 : begin
        result = input_748;
      end
      11'b01011101101 : begin
        result = input_749;
      end
      11'b01011101110 : begin
        result = input_750;
      end
      11'b01011101111 : begin
        result = input_751;
      end
      11'b01011110000 : begin
        result = input_752;
      end
      11'b01011110001 : begin
        result = input_753;
      end
      11'b01011110010 : begin
        result = input_754;
      end
      11'b01011110011 : begin
        result = input_755;
      end
      11'b01011110100 : begin
        result = input_756;
      end
      11'b01011110101 : begin
        result = input_757;
      end
      11'b01011110110 : begin
        result = input_758;
      end
      11'b01011110111 : begin
        result = input_759;
      end
      11'b01011111000 : begin
        result = input_760;
      end
      11'b01011111001 : begin
        result = input_761;
      end
      11'b01011111010 : begin
        result = input_762;
      end
      11'b01011111011 : begin
        result = input_763;
      end
      11'b01011111100 : begin
        result = input_764;
      end
      11'b01011111101 : begin
        result = input_765;
      end
      11'b01011111110 : begin
        result = input_766;
      end
      11'b01011111111 : begin
        result = input_767;
      end
      11'b01100000000 : begin
        result = input_768;
      end
      11'b01100000001 : begin
        result = input_769;
      end
      11'b01100000010 : begin
        result = input_770;
      end
      11'b01100000011 : begin
        result = input_771;
      end
      11'b01100000100 : begin
        result = input_772;
      end
      11'b01100000101 : begin
        result = input_773;
      end
      11'b01100000110 : begin
        result = input_774;
      end
      11'b01100000111 : begin
        result = input_775;
      end
      11'b01100001000 : begin
        result = input_776;
      end
      11'b01100001001 : begin
        result = input_777;
      end
      11'b01100001010 : begin
        result = input_778;
      end
      11'b01100001011 : begin
        result = input_779;
      end
      11'b01100001100 : begin
        result = input_780;
      end
      11'b01100001101 : begin
        result = input_781;
      end
      11'b01100001110 : begin
        result = input_782;
      end
      11'b01100001111 : begin
        result = input_783;
      end
      11'b01100010000 : begin
        result = input_784;
      end
      11'b01100010001 : begin
        result = input_785;
      end
      11'b01100010010 : begin
        result = input_786;
      end
      11'b01100010011 : begin
        result = input_787;
      end
      11'b01100010100 : begin
        result = input_788;
      end
      11'b01100010101 : begin
        result = input_789;
      end
      11'b01100010110 : begin
        result = input_790;
      end
      11'b01100010111 : begin
        result = input_791;
      end
      11'b01100011000 : begin
        result = input_792;
      end
      11'b01100011001 : begin
        result = input_793;
      end
      11'b01100011010 : begin
        result = input_794;
      end
      11'b01100011011 : begin
        result = input_795;
      end
      11'b01100011100 : begin
        result = input_796;
      end
      11'b01100011101 : begin
        result = input_797;
      end
      11'b01100011110 : begin
        result = input_798;
      end
      11'b01100011111 : begin
        result = input_799;
      end
      11'b01100100000 : begin
        result = input_800;
      end
      11'b01100100001 : begin
        result = input_801;
      end
      11'b01100100010 : begin
        result = input_802;
      end
      11'b01100100011 : begin
        result = input_803;
      end
      11'b01100100100 : begin
        result = input_804;
      end
      11'b01100100101 : begin
        result = input_805;
      end
      11'b01100100110 : begin
        result = input_806;
      end
      11'b01100100111 : begin
        result = input_807;
      end
      11'b01100101000 : begin
        result = input_808;
      end
      11'b01100101001 : begin
        result = input_809;
      end
      11'b01100101010 : begin
        result = input_810;
      end
      11'b01100101011 : begin
        result = input_811;
      end
      11'b01100101100 : begin
        result = input_812;
      end
      11'b01100101101 : begin
        result = input_813;
      end
      11'b01100101110 : begin
        result = input_814;
      end
      11'b01100101111 : begin
        result = input_815;
      end
      11'b01100110000 : begin
        result = input_816;
      end
      11'b01100110001 : begin
        result = input_817;
      end
      11'b01100110010 : begin
        result = input_818;
      end
      11'b01100110011 : begin
        result = input_819;
      end
      11'b01100110100 : begin
        result = input_820;
      end
      11'b01100110101 : begin
        result = input_821;
      end
      11'b01100110110 : begin
        result = input_822;
      end
      11'b01100110111 : begin
        result = input_823;
      end
      11'b01100111000 : begin
        result = input_824;
      end
      11'b01100111001 : begin
        result = input_825;
      end
      11'b01100111010 : begin
        result = input_826;
      end
      11'b01100111011 : begin
        result = input_827;
      end
      11'b01100111100 : begin
        result = input_828;
      end
      11'b01100111101 : begin
        result = input_829;
      end
      11'b01100111110 : begin
        result = input_830;
      end
      11'b01100111111 : begin
        result = input_831;
      end
      11'b01101000000 : begin
        result = input_832;
      end
      11'b01101000001 : begin
        result = input_833;
      end
      11'b01101000010 : begin
        result = input_834;
      end
      11'b01101000011 : begin
        result = input_835;
      end
      11'b01101000100 : begin
        result = input_836;
      end
      11'b01101000101 : begin
        result = input_837;
      end
      11'b01101000110 : begin
        result = input_838;
      end
      11'b01101000111 : begin
        result = input_839;
      end
      11'b01101001000 : begin
        result = input_840;
      end
      11'b01101001001 : begin
        result = input_841;
      end
      11'b01101001010 : begin
        result = input_842;
      end
      11'b01101001011 : begin
        result = input_843;
      end
      11'b01101001100 : begin
        result = input_844;
      end
      11'b01101001101 : begin
        result = input_845;
      end
      11'b01101001110 : begin
        result = input_846;
      end
      11'b01101001111 : begin
        result = input_847;
      end
      11'b01101010000 : begin
        result = input_848;
      end
      11'b01101010001 : begin
        result = input_849;
      end
      11'b01101010010 : begin
        result = input_850;
      end
      11'b01101010011 : begin
        result = input_851;
      end
      11'b01101010100 : begin
        result = input_852;
      end
      11'b01101010101 : begin
        result = input_853;
      end
      11'b01101010110 : begin
        result = input_854;
      end
      11'b01101010111 : begin
        result = input_855;
      end
      11'b01101011000 : begin
        result = input_856;
      end
      11'b01101011001 : begin
        result = input_857;
      end
      11'b01101011010 : begin
        result = input_858;
      end
      11'b01101011011 : begin
        result = input_859;
      end
      11'b01101011100 : begin
        result = input_860;
      end
      11'b01101011101 : begin
        result = input_861;
      end
      11'b01101011110 : begin
        result = input_862;
      end
      11'b01101011111 : begin
        result = input_863;
      end
      11'b01101100000 : begin
        result = input_864;
      end
      11'b01101100001 : begin
        result = input_865;
      end
      11'b01101100010 : begin
        result = input_866;
      end
      11'b01101100011 : begin
        result = input_867;
      end
      11'b01101100100 : begin
        result = input_868;
      end
      11'b01101100101 : begin
        result = input_869;
      end
      11'b01101100110 : begin
        result = input_870;
      end
      11'b01101100111 : begin
        result = input_871;
      end
      11'b01101101000 : begin
        result = input_872;
      end
      11'b01101101001 : begin
        result = input_873;
      end
      11'b01101101010 : begin
        result = input_874;
      end
      11'b01101101011 : begin
        result = input_875;
      end
      11'b01101101100 : begin
        result = input_876;
      end
      11'b01101101101 : begin
        result = input_877;
      end
      11'b01101101110 : begin
        result = input_878;
      end
      11'b01101101111 : begin
        result = input_879;
      end
      11'b01101110000 : begin
        result = input_880;
      end
      11'b01101110001 : begin
        result = input_881;
      end
      11'b01101110010 : begin
        result = input_882;
      end
      11'b01101110011 : begin
        result = input_883;
      end
      11'b01101110100 : begin
        result = input_884;
      end
      11'b01101110101 : begin
        result = input_885;
      end
      11'b01101110110 : begin
        result = input_886;
      end
      11'b01101110111 : begin
        result = input_887;
      end
      11'b01101111000 : begin
        result = input_888;
      end
      11'b01101111001 : begin
        result = input_889;
      end
      11'b01101111010 : begin
        result = input_890;
      end
      11'b01101111011 : begin
        result = input_891;
      end
      11'b01101111100 : begin
        result = input_892;
      end
      11'b01101111101 : begin
        result = input_893;
      end
      11'b01101111110 : begin
        result = input_894;
      end
      11'b01101111111 : begin
        result = input_895;
      end
      11'b01110000000 : begin
        result = input_896;
      end
      11'b01110000001 : begin
        result = input_897;
      end
      11'b01110000010 : begin
        result = input_898;
      end
      11'b01110000011 : begin
        result = input_899;
      end
      11'b01110000100 : begin
        result = input_900;
      end
      11'b01110000101 : begin
        result = input_901;
      end
      11'b01110000110 : begin
        result = input_902;
      end
      11'b01110000111 : begin
        result = input_903;
      end
      11'b01110001000 : begin
        result = input_904;
      end
      11'b01110001001 : begin
        result = input_905;
      end
      11'b01110001010 : begin
        result = input_906;
      end
      11'b01110001011 : begin
        result = input_907;
      end
      11'b01110001100 : begin
        result = input_908;
      end
      11'b01110001101 : begin
        result = input_909;
      end
      11'b01110001110 : begin
        result = input_910;
      end
      11'b01110001111 : begin
        result = input_911;
      end
      11'b01110010000 : begin
        result = input_912;
      end
      11'b01110010001 : begin
        result = input_913;
      end
      11'b01110010010 : begin
        result = input_914;
      end
      11'b01110010011 : begin
        result = input_915;
      end
      11'b01110010100 : begin
        result = input_916;
      end
      11'b01110010101 : begin
        result = input_917;
      end
      11'b01110010110 : begin
        result = input_918;
      end
      11'b01110010111 : begin
        result = input_919;
      end
      11'b01110011000 : begin
        result = input_920;
      end
      11'b01110011001 : begin
        result = input_921;
      end
      11'b01110011010 : begin
        result = input_922;
      end
      11'b01110011011 : begin
        result = input_923;
      end
      11'b01110011100 : begin
        result = input_924;
      end
      11'b01110011101 : begin
        result = input_925;
      end
      11'b01110011110 : begin
        result = input_926;
      end
      11'b01110011111 : begin
        result = input_927;
      end
      11'b01110100000 : begin
        result = input_928;
      end
      11'b01110100001 : begin
        result = input_929;
      end
      11'b01110100010 : begin
        result = input_930;
      end
      11'b01110100011 : begin
        result = input_931;
      end
      11'b01110100100 : begin
        result = input_932;
      end
      11'b01110100101 : begin
        result = input_933;
      end
      11'b01110100110 : begin
        result = input_934;
      end
      11'b01110100111 : begin
        result = input_935;
      end
      11'b01110101000 : begin
        result = input_936;
      end
      11'b01110101001 : begin
        result = input_937;
      end
      11'b01110101010 : begin
        result = input_938;
      end
      11'b01110101011 : begin
        result = input_939;
      end
      11'b01110101100 : begin
        result = input_940;
      end
      11'b01110101101 : begin
        result = input_941;
      end
      11'b01110101110 : begin
        result = input_942;
      end
      11'b01110101111 : begin
        result = input_943;
      end
      11'b01110110000 : begin
        result = input_944;
      end
      11'b01110110001 : begin
        result = input_945;
      end
      11'b01110110010 : begin
        result = input_946;
      end
      11'b01110110011 : begin
        result = input_947;
      end
      11'b01110110100 : begin
        result = input_948;
      end
      11'b01110110101 : begin
        result = input_949;
      end
      11'b01110110110 : begin
        result = input_950;
      end
      11'b01110110111 : begin
        result = input_951;
      end
      11'b01110111000 : begin
        result = input_952;
      end
      11'b01110111001 : begin
        result = input_953;
      end
      11'b01110111010 : begin
        result = input_954;
      end
      11'b01110111011 : begin
        result = input_955;
      end
      11'b01110111100 : begin
        result = input_956;
      end
      11'b01110111101 : begin
        result = input_957;
      end
      11'b01110111110 : begin
        result = input_958;
      end
      11'b01110111111 : begin
        result = input_959;
      end
      11'b01111000000 : begin
        result = input_960;
      end
      11'b01111000001 : begin
        result = input_961;
      end
      11'b01111000010 : begin
        result = input_962;
      end
      11'b01111000011 : begin
        result = input_963;
      end
      11'b01111000100 : begin
        result = input_964;
      end
      11'b01111000101 : begin
        result = input_965;
      end
      11'b01111000110 : begin
        result = input_966;
      end
      11'b01111000111 : begin
        result = input_967;
      end
      11'b01111001000 : begin
        result = input_968;
      end
      11'b01111001001 : begin
        result = input_969;
      end
      11'b01111001010 : begin
        result = input_970;
      end
      11'b01111001011 : begin
        result = input_971;
      end
      11'b01111001100 : begin
        result = input_972;
      end
      11'b01111001101 : begin
        result = input_973;
      end
      11'b01111001110 : begin
        result = input_974;
      end
      11'b01111001111 : begin
        result = input_975;
      end
      11'b01111010000 : begin
        result = input_976;
      end
      11'b01111010001 : begin
        result = input_977;
      end
      11'b01111010010 : begin
        result = input_978;
      end
      11'b01111010011 : begin
        result = input_979;
      end
      11'b01111010100 : begin
        result = input_980;
      end
      11'b01111010101 : begin
        result = input_981;
      end
      11'b01111010110 : begin
        result = input_982;
      end
      11'b01111010111 : begin
        result = input_983;
      end
      11'b01111011000 : begin
        result = input_984;
      end
      11'b01111011001 : begin
        result = input_985;
      end
      11'b01111011010 : begin
        result = input_986;
      end
      11'b01111011011 : begin
        result = input_987;
      end
      11'b01111011100 : begin
        result = input_988;
      end
      11'b01111011101 : begin
        result = input_989;
      end
      11'b01111011110 : begin
        result = input_990;
      end
      11'b01111011111 : begin
        result = input_991;
      end
      11'b01111100000 : begin
        result = input_992;
      end
      11'b01111100001 : begin
        result = input_993;
      end
      11'b01111100010 : begin
        result = input_994;
      end
      11'b01111100011 : begin
        result = input_995;
      end
      11'b01111100100 : begin
        result = input_996;
      end
      11'b01111100101 : begin
        result = input_997;
      end
      11'b01111100110 : begin
        result = input_998;
      end
      11'b01111100111 : begin
        result = input_999;
      end
      11'b01111101000 : begin
        result = input_1000;
      end
      11'b01111101001 : begin
        result = input_1001;
      end
      11'b01111101010 : begin
        result = input_1002;
      end
      11'b01111101011 : begin
        result = input_1003;
      end
      11'b01111101100 : begin
        result = input_1004;
      end
      11'b01111101101 : begin
        result = input_1005;
      end
      11'b01111101110 : begin
        result = input_1006;
      end
      11'b01111101111 : begin
        result = input_1007;
      end
      11'b01111110000 : begin
        result = input_1008;
      end
      11'b01111110001 : begin
        result = input_1009;
      end
      11'b01111110010 : begin
        result = input_1010;
      end
      11'b01111110011 : begin
        result = input_1011;
      end
      11'b01111110100 : begin
        result = input_1012;
      end
      11'b01111110101 : begin
        result = input_1013;
      end
      11'b01111110110 : begin
        result = input_1014;
      end
      11'b01111110111 : begin
        result = input_1015;
      end
      11'b01111111000 : begin
        result = input_1016;
      end
      11'b01111111001 : begin
        result = input_1017;
      end
      11'b01111111010 : begin
        result = input_1018;
      end
      11'b01111111011 : begin
        result = input_1019;
      end
      11'b01111111100 : begin
        result = input_1020;
      end
      11'b01111111101 : begin
        result = input_1021;
      end
      11'b01111111110 : begin
        result = input_1022;
      end
      11'b01111111111 : begin
        result = input_1023;
      end
      11'b10000000000 : begin
        result = input_1024;
      end
      11'b10000000001 : begin
        result = input_1025;
      end
      11'b10000000010 : begin
        result = input_1026;
      end
      11'b10000000011 : begin
        result = input_1027;
      end
      11'b10000000100 : begin
        result = input_1028;
      end
      11'b10000000101 : begin
        result = input_1029;
      end
      11'b10000000110 : begin
        result = input_1030;
      end
      11'b10000000111 : begin
        result = input_1031;
      end
      11'b10000001000 : begin
        result = input_1032;
      end
      11'b10000001001 : begin
        result = input_1033;
      end
      11'b10000001010 : begin
        result = input_1034;
      end
      11'b10000001011 : begin
        result = input_1035;
      end
      11'b10000001100 : begin
        result = input_1036;
      end
      11'b10000001101 : begin
        result = input_1037;
      end
      11'b10000001110 : begin
        result = input_1038;
      end
      11'b10000001111 : begin
        result = input_1039;
      end
      11'b10000010000 : begin
        result = input_1040;
      end
      11'b10000010001 : begin
        result = input_1041;
      end
      11'b10000010010 : begin
        result = input_1042;
      end
      11'b10000010011 : begin
        result = input_1043;
      end
      11'b10000010100 : begin
        result = input_1044;
      end
      11'b10000010101 : begin
        result = input_1045;
      end
      11'b10000010110 : begin
        result = input_1046;
      end
      11'b10000010111 : begin
        result = input_1047;
      end
      11'b10000011000 : begin
        result = input_1048;
      end
      11'b10000011001 : begin
        result = input_1049;
      end
      11'b10000011010 : begin
        result = input_1050;
      end
      11'b10000011011 : begin
        result = input_1051;
      end
      11'b10000011100 : begin
        result = input_1052;
      end
      11'b10000011101 : begin
        result = input_1053;
      end
      11'b10000011110 : begin
        result = input_1054;
      end
      11'b10000011111 : begin
        result = input_1055;
      end
      11'b10000100000 : begin
        result = input_1056;
      end
      11'b10000100001 : begin
        result = input_1057;
      end
      11'b10000100010 : begin
        result = input_1058;
      end
      11'b10000100011 : begin
        result = input_1059;
      end
      11'b10000100100 : begin
        result = input_1060;
      end
      11'b10000100101 : begin
        result = input_1061;
      end
      11'b10000100110 : begin
        result = input_1062;
      end
      11'b10000100111 : begin
        result = input_1063;
      end
      11'b10000101000 : begin
        result = input_1064;
      end
      11'b10000101001 : begin
        result = input_1065;
      end
      11'b10000101010 : begin
        result = input_1066;
      end
      11'b10000101011 : begin
        result = input_1067;
      end
      11'b10000101100 : begin
        result = input_1068;
      end
      11'b10000101101 : begin
        result = input_1069;
      end
      11'b10000101110 : begin
        result = input_1070;
      end
      11'b10000101111 : begin
        result = input_1071;
      end
      11'b10000110000 : begin
        result = input_1072;
      end
      11'b10000110001 : begin
        result = input_1073;
      end
      11'b10000110010 : begin
        result = input_1074;
      end
      11'b10000110011 : begin
        result = input_1075;
      end
      11'b10000110100 : begin
        result = input_1076;
      end
      11'b10000110101 : begin
        result = input_1077;
      end
      11'b10000110110 : begin
        result = input_1078;
      end
      11'b10000110111 : begin
        result = input_1079;
      end
      11'b10000111000 : begin
        result = input_1080;
      end
      11'b10000111001 : begin
        result = input_1081;
      end
      11'b10000111010 : begin
        result = input_1082;
      end
      11'b10000111011 : begin
        result = input_1083;
      end
      11'b10000111100 : begin
        result = input_1084;
      end
      11'b10000111101 : begin
        result = input_1085;
      end
      11'b10000111110 : begin
        result = input_1086;
      end
      11'b10000111111 : begin
        result = input_1087;
      end
      11'b10001000000 : begin
        result = input_1088;
      end
      11'b10001000001 : begin
        result = input_1089;
      end
      11'b10001000010 : begin
        result = input_1090;
      end
      11'b10001000011 : begin
        result = input_1091;
      end
      11'b10001000100 : begin
        result = input_1092;
      end
      11'b10001000101 : begin
        result = input_1093;
      end
      11'b10001000110 : begin
        result = input_1094;
      end
      11'b10001000111 : begin
        result = input_1095;
      end
      11'b10001001000 : begin
        result = input_1096;
      end
      11'b10001001001 : begin
        result = input_1097;
      end
      11'b10001001010 : begin
        result = input_1098;
      end
      11'b10001001011 : begin
        result = input_1099;
      end
      11'b10001001100 : begin
        result = input_1100;
      end
      11'b10001001101 : begin
        result = input_1101;
      end
      11'b10001001110 : begin
        result = input_1102;
      end
      11'b10001001111 : begin
        result = input_1103;
      end
      11'b10001010000 : begin
        result = input_1104;
      end
      11'b10001010001 : begin
        result = input_1105;
      end
      11'b10001010010 : begin
        result = input_1106;
      end
      11'b10001010011 : begin
        result = input_1107;
      end
      11'b10001010100 : begin
        result = input_1108;
      end
      11'b10001010101 : begin
        result = input_1109;
      end
      11'b10001010110 : begin
        result = input_1110;
      end
      11'b10001010111 : begin
        result = input_1111;
      end
      11'b10001011000 : begin
        result = input_1112;
      end
      11'b10001011001 : begin
        result = input_1113;
      end
      11'b10001011010 : begin
        result = input_1114;
      end
      11'b10001011011 : begin
        result = input_1115;
      end
      11'b10001011100 : begin
        result = input_1116;
      end
      11'b10001011101 : begin
        result = input_1117;
      end
      11'b10001011110 : begin
        result = input_1118;
      end
      11'b10001011111 : begin
        result = input_1119;
      end
      11'b10001100000 : begin
        result = input_1120;
      end
      11'b10001100001 : begin
        result = input_1121;
      end
      11'b10001100010 : begin
        result = input_1122;
      end
      11'b10001100011 : begin
        result = input_1123;
      end
      11'b10001100100 : begin
        result = input_1124;
      end
      11'b10001100101 : begin
        result = input_1125;
      end
      11'b10001100110 : begin
        result = input_1126;
      end
      11'b10001100111 : begin
        result = input_1127;
      end
      11'b10001101000 : begin
        result = input_1128;
      end
      11'b10001101001 : begin
        result = input_1129;
      end
      11'b10001101010 : begin
        result = input_1130;
      end
      11'b10001101011 : begin
        result = input_1131;
      end
      11'b10001101100 : begin
        result = input_1132;
      end
      11'b10001101101 : begin
        result = input_1133;
      end
      11'b10001101110 : begin
        result = input_1134;
      end
      11'b10001101111 : begin
        result = input_1135;
      end
      11'b10001110000 : begin
        result = input_1136;
      end
      11'b10001110001 : begin
        result = input_1137;
      end
      11'b10001110010 : begin
        result = input_1138;
      end
      11'b10001110011 : begin
        result = input_1139;
      end
      11'b10001110100 : begin
        result = input_1140;
      end
      11'b10001110101 : begin
        result = input_1141;
      end
      11'b10001110110 : begin
        result = input_1142;
      end
      11'b10001110111 : begin
        result = input_1143;
      end
      11'b10001111000 : begin
        result = input_1144;
      end
      11'b10001111001 : begin
        result = input_1145;
      end
      11'b10001111010 : begin
        result = input_1146;
      end
      11'b10001111011 : begin
        result = input_1147;
      end
      11'b10001111100 : begin
        result = input_1148;
      end
      11'b10001111101 : begin
        result = input_1149;
      end
      11'b10001111110 : begin
        result = input_1150;
      end
      11'b10001111111 : begin
        result = input_1151;
      end
      11'b10010000000 : begin
        result = input_1152;
      end
      11'b10010000001 : begin
        result = input_1153;
      end
      11'b10010000010 : begin
        result = input_1154;
      end
      11'b10010000011 : begin
        result = input_1155;
      end
      11'b10010000100 : begin
        result = input_1156;
      end
      11'b10010000101 : begin
        result = input_1157;
      end
      11'b10010000110 : begin
        result = input_1158;
      end
      11'b10010000111 : begin
        result = input_1159;
      end
      11'b10010001000 : begin
        result = input_1160;
      end
      11'b10010001001 : begin
        result = input_1161;
      end
      11'b10010001010 : begin
        result = input_1162;
      end
      11'b10010001011 : begin
        result = input_1163;
      end
      11'b10010001100 : begin
        result = input_1164;
      end
      11'b10010001101 : begin
        result = input_1165;
      end
      11'b10010001110 : begin
        result = input_1166;
      end
      11'b10010001111 : begin
        result = input_1167;
      end
      11'b10010010000 : begin
        result = input_1168;
      end
      11'b10010010001 : begin
        result = input_1169;
      end
      11'b10010010010 : begin
        result = input_1170;
      end
      11'b10010010011 : begin
        result = input_1171;
      end
      11'b10010010100 : begin
        result = input_1172;
      end
      11'b10010010101 : begin
        result = input_1173;
      end
      11'b10010010110 : begin
        result = input_1174;
      end
      11'b10010010111 : begin
        result = input_1175;
      end
      11'b10010011000 : begin
        result = input_1176;
      end
      11'b10010011001 : begin
        result = input_1177;
      end
      11'b10010011010 : begin
        result = input_1178;
      end
      11'b10010011011 : begin
        result = input_1179;
      end
      11'b10010011100 : begin
        result = input_1180;
      end
      11'b10010011101 : begin
        result = input_1181;
      end
      11'b10010011110 : begin
        result = input_1182;
      end
      11'b10010011111 : begin
        result = input_1183;
      end
      11'b10010100000 : begin
        result = input_1184;
      end
      11'b10010100001 : begin
        result = input_1185;
      end
      11'b10010100010 : begin
        result = input_1186;
      end
      11'b10010100011 : begin
        result = input_1187;
      end
      11'b10010100100 : begin
        result = input_1188;
      end
      11'b10010100101 : begin
        result = input_1189;
      end
      11'b10010100110 : begin
        result = input_1190;
      end
      11'b10010100111 : begin
        result = input_1191;
      end
      11'b10010101000 : begin
        result = input_1192;
      end
      11'b10010101001 : begin
        result = input_1193;
      end
      11'b10010101010 : begin
        result = input_1194;
      end
      11'b10010101011 : begin
        result = input_1195;
      end
      11'b10010101100 : begin
        result = input_1196;
      end
      11'b10010101101 : begin
        result = input_1197;
      end
      11'b10010101110 : begin
        result = input_1198;
      end
      11'b10010101111 : begin
        result = input_1199;
      end
      11'b10010110000 : begin
        result = input_1200;
      end
      11'b10010110001 : begin
        result = input_1201;
      end
      11'b10010110010 : begin
        result = input_1202;
      end
      11'b10010110011 : begin
        result = input_1203;
      end
      11'b10010110100 : begin
        result = input_1204;
      end
      11'b10010110101 : begin
        result = input_1205;
      end
      11'b10010110110 : begin
        result = input_1206;
      end
      11'b10010110111 : begin
        result = input_1207;
      end
      11'b10010111000 : begin
        result = input_1208;
      end
      11'b10010111001 : begin
        result = input_1209;
      end
      11'b10010111010 : begin
        result = input_1210;
      end
      11'b10010111011 : begin
        result = input_1211;
      end
      11'b10010111100 : begin
        result = input_1212;
      end
      11'b10010111101 : begin
        result = input_1213;
      end
      11'b10010111110 : begin
        result = input_1214;
      end
      11'b10010111111 : begin
        result = input_1215;
      end
      11'b10011000000 : begin
        result = input_1216;
      end
      11'b10011000001 : begin
        result = input_1217;
      end
      11'b10011000010 : begin
        result = input_1218;
      end
      11'b10011000011 : begin
        result = input_1219;
      end
      11'b10011000100 : begin
        result = input_1220;
      end
      11'b10011000101 : begin
        result = input_1221;
      end
      11'b10011000110 : begin
        result = input_1222;
      end
      11'b10011000111 : begin
        result = input_1223;
      end
      11'b10011001000 : begin
        result = input_1224;
      end
      11'b10011001001 : begin
        result = input_1225;
      end
      11'b10011001010 : begin
        result = input_1226;
      end
      11'b10011001011 : begin
        result = input_1227;
      end
      11'b10011001100 : begin
        result = input_1228;
      end
      11'b10011001101 : begin
        result = input_1229;
      end
      11'b10011001110 : begin
        result = input_1230;
      end
      11'b10011001111 : begin
        result = input_1231;
      end
      11'b10011010000 : begin
        result = input_1232;
      end
      11'b10011010001 : begin
        result = input_1233;
      end
      11'b10011010010 : begin
        result = input_1234;
      end
      11'b10011010011 : begin
        result = input_1235;
      end
      11'b10011010100 : begin
        result = input_1236;
      end
      11'b10011010101 : begin
        result = input_1237;
      end
      11'b10011010110 : begin
        result = input_1238;
      end
      11'b10011010111 : begin
        result = input_1239;
      end
      11'b10011011000 : begin
        result = input_1240;
      end
      11'b10011011001 : begin
        result = input_1241;
      end
      11'b10011011010 : begin
        result = input_1242;
      end
      11'b10011011011 : begin
        result = input_1243;
      end
      11'b10011011100 : begin
        result = input_1244;
      end
      11'b10011011101 : begin
        result = input_1245;
      end
      11'b10011011110 : begin
        result = input_1246;
      end
      11'b10011011111 : begin
        result = input_1247;
      end
      11'b10011100000 : begin
        result = input_1248;
      end
      11'b10011100001 : begin
        result = input_1249;
      end
      11'b10011100010 : begin
        result = input_1250;
      end
      11'b10011100011 : begin
        result = input_1251;
      end
      11'b10011100100 : begin
        result = input_1252;
      end
      11'b10011100101 : begin
        result = input_1253;
      end
      11'b10011100110 : begin
        result = input_1254;
      end
      11'b10011100111 : begin
        result = input_1255;
      end
      11'b10011101000 : begin
        result = input_1256;
      end
      11'b10011101001 : begin
        result = input_1257;
      end
      11'b10011101010 : begin
        result = input_1258;
      end
      11'b10011101011 : begin
        result = input_1259;
      end
      11'b10011101100 : begin
        result = input_1260;
      end
      11'b10011101101 : begin
        result = input_1261;
      end
      11'b10011101110 : begin
        result = input_1262;
      end
      11'b10011101111 : begin
        result = input_1263;
      end
      11'b10011110000 : begin
        result = input_1264;
      end
      11'b10011110001 : begin
        result = input_1265;
      end
      11'b10011110010 : begin
        result = input_1266;
      end
      11'b10011110011 : begin
        result = input_1267;
      end
      11'b10011110100 : begin
        result = input_1268;
      end
      11'b10011110101 : begin
        result = input_1269;
      end
      11'b10011110110 : begin
        result = input_1270;
      end
      11'b10011110111 : begin
        result = input_1271;
      end
      11'b10011111000 : begin
        result = input_1272;
      end
      11'b10011111001 : begin
        result = input_1273;
      end
      11'b10011111010 : begin
        result = input_1274;
      end
      11'b10011111011 : begin
        result = input_1275;
      end
      11'b10011111100 : begin
        result = input_1276;
      end
      11'b10011111101 : begin
        result = input_1277;
      end
      11'b10011111110 : begin
        result = input_1278;
      end
      11'b10011111111 : begin
        result = input_1279;
      end
      11'b10100000000 : begin
        result = input_1280;
      end
      11'b10100000001 : begin
        result = input_1281;
      end
      11'b10100000010 : begin
        result = input_1282;
      end
      11'b10100000011 : begin
        result = input_1283;
      end
      11'b10100000100 : begin
        result = input_1284;
      end
      11'b10100000101 : begin
        result = input_1285;
      end
      11'b10100000110 : begin
        result = input_1286;
      end
      11'b10100000111 : begin
        result = input_1287;
      end
      11'b10100001000 : begin
        result = input_1288;
      end
      11'b10100001001 : begin
        result = input_1289;
      end
      11'b10100001010 : begin
        result = input_1290;
      end
      11'b10100001011 : begin
        result = input_1291;
      end
      11'b10100001100 : begin
        result = input_1292;
      end
      11'b10100001101 : begin
        result = input_1293;
      end
      11'b10100001110 : begin
        result = input_1294;
      end
      11'b10100001111 : begin
        result = input_1295;
      end
      11'b10100010000 : begin
        result = input_1296;
      end
      11'b10100010001 : begin
        result = input_1297;
      end
      11'b10100010010 : begin
        result = input_1298;
      end
      11'b10100010011 : begin
        result = input_1299;
      end
      11'b10100010100 : begin
        result = input_1300;
      end
      11'b10100010101 : begin
        result = input_1301;
      end
      11'b10100010110 : begin
        result = input_1302;
      end
      11'b10100010111 : begin
        result = input_1303;
      end
      11'b10100011000 : begin
        result = input_1304;
      end
      11'b10100011001 : begin
        result = input_1305;
      end
      11'b10100011010 : begin
        result = input_1306;
      end
      11'b10100011011 : begin
        result = input_1307;
      end
      11'b10100011100 : begin
        result = input_1308;
      end
      11'b10100011101 : begin
        result = input_1309;
      end
      11'b10100011110 : begin
        result = input_1310;
      end
      11'b10100011111 : begin
        result = input_1311;
      end
      11'b10100100000 : begin
        result = input_1312;
      end
      11'b10100100001 : begin
        result = input_1313;
      end
      11'b10100100010 : begin
        result = input_1314;
      end
      11'b10100100011 : begin
        result = input_1315;
      end
      11'b10100100100 : begin
        result = input_1316;
      end
      11'b10100100101 : begin
        result = input_1317;
      end
      11'b10100100110 : begin
        result = input_1318;
      end
      11'b10100100111 : begin
        result = input_1319;
      end
      11'b10100101000 : begin
        result = input_1320;
      end
      11'b10100101001 : begin
        result = input_1321;
      end
      11'b10100101010 : begin
        result = input_1322;
      end
      11'b10100101011 : begin
        result = input_1323;
      end
      11'b10100101100 : begin
        result = input_1324;
      end
      11'b10100101101 : begin
        result = input_1325;
      end
      11'b10100101110 : begin
        result = input_1326;
      end
      11'b10100101111 : begin
        result = input_1327;
      end
      11'b10100110000 : begin
        result = input_1328;
      end
      11'b10100110001 : begin
        result = input_1329;
      end
      11'b10100110010 : begin
        result = input_1330;
      end
      11'b10100110011 : begin
        result = input_1331;
      end
      11'b10100110100 : begin
        result = input_1332;
      end
      11'b10100110101 : begin
        result = input_1333;
      end
      11'b10100110110 : begin
        result = input_1334;
      end
      11'b10100110111 : begin
        result = input_1335;
      end
      11'b10100111000 : begin
        result = input_1336;
      end
      11'b10100111001 : begin
        result = input_1337;
      end
      11'b10100111010 : begin
        result = input_1338;
      end
      11'b10100111011 : begin
        result = input_1339;
      end
      11'b10100111100 : begin
        result = input_1340;
      end
      11'b10100111101 : begin
        result = input_1341;
      end
      11'b10100111110 : begin
        result = input_1342;
      end
      11'b10100111111 : begin
        result = input_1343;
      end
      11'b10101000000 : begin
        result = input_1344;
      end
      11'b10101000001 : begin
        result = input_1345;
      end
      11'b10101000010 : begin
        result = input_1346;
      end
      11'b10101000011 : begin
        result = input_1347;
      end
      11'b10101000100 : begin
        result = input_1348;
      end
      11'b10101000101 : begin
        result = input_1349;
      end
      11'b10101000110 : begin
        result = input_1350;
      end
      11'b10101000111 : begin
        result = input_1351;
      end
      11'b10101001000 : begin
        result = input_1352;
      end
      11'b10101001001 : begin
        result = input_1353;
      end
      11'b10101001010 : begin
        result = input_1354;
      end
      11'b10101001011 : begin
        result = input_1355;
      end
      11'b10101001100 : begin
        result = input_1356;
      end
      11'b10101001101 : begin
        result = input_1357;
      end
      11'b10101001110 : begin
        result = input_1358;
      end
      11'b10101001111 : begin
        result = input_1359;
      end
      11'b10101010000 : begin
        result = input_1360;
      end
      11'b10101010001 : begin
        result = input_1361;
      end
      11'b10101010010 : begin
        result = input_1362;
      end
      11'b10101010011 : begin
        result = input_1363;
      end
      11'b10101010100 : begin
        result = input_1364;
      end
      11'b10101010101 : begin
        result = input_1365;
      end
      11'b10101010110 : begin
        result = input_1366;
      end
      11'b10101010111 : begin
        result = input_1367;
      end
      11'b10101011000 : begin
        result = input_1368;
      end
      11'b10101011001 : begin
        result = input_1369;
      end
      11'b10101011010 : begin
        result = input_1370;
      end
      11'b10101011011 : begin
        result = input_1371;
      end
      11'b10101011100 : begin
        result = input_1372;
      end
      11'b10101011101 : begin
        result = input_1373;
      end
      11'b10101011110 : begin
        result = input_1374;
      end
      11'b10101011111 : begin
        result = input_1375;
      end
      11'b10101100000 : begin
        result = input_1376;
      end
      11'b10101100001 : begin
        result = input_1377;
      end
      11'b10101100010 : begin
        result = input_1378;
      end
      11'b10101100011 : begin
        result = input_1379;
      end
      11'b10101100100 : begin
        result = input_1380;
      end
      11'b10101100101 : begin
        result = input_1381;
      end
      11'b10101100110 : begin
        result = input_1382;
      end
      11'b10101100111 : begin
        result = input_1383;
      end
      11'b10101101000 : begin
        result = input_1384;
      end
      11'b10101101001 : begin
        result = input_1385;
      end
      11'b10101101010 : begin
        result = input_1386;
      end
      11'b10101101011 : begin
        result = input_1387;
      end
      11'b10101101100 : begin
        result = input_1388;
      end
      11'b10101101101 : begin
        result = input_1389;
      end
      11'b10101101110 : begin
        result = input_1390;
      end
      11'b10101101111 : begin
        result = input_1391;
      end
      11'b10101110000 : begin
        result = input_1392;
      end
      11'b10101110001 : begin
        result = input_1393;
      end
      11'b10101110010 : begin
        result = input_1394;
      end
      11'b10101110011 : begin
        result = input_1395;
      end
      11'b10101110100 : begin
        result = input_1396;
      end
      11'b10101110101 : begin
        result = input_1397;
      end
      11'b10101110110 : begin
        result = input_1398;
      end
      11'b10101110111 : begin
        result = input_1399;
      end
      11'b10101111000 : begin
        result = input_1400;
      end
      11'b10101111001 : begin
        result = input_1401;
      end
      11'b10101111010 : begin
        result = input_1402;
      end
      11'b10101111011 : begin
        result = input_1403;
      end
      11'b10101111100 : begin
        result = input_1404;
      end
      11'b10101111101 : begin
        result = input_1405;
      end
      11'b10101111110 : begin
        result = input_1406;
      end
      11'b10101111111 : begin
        result = input_1407;
      end
      11'b10110000000 : begin
        result = input_1408;
      end
      11'b10110000001 : begin
        result = input_1409;
      end
      11'b10110000010 : begin
        result = input_1410;
      end
      11'b10110000011 : begin
        result = input_1411;
      end
      11'b10110000100 : begin
        result = input_1412;
      end
      11'b10110000101 : begin
        result = input_1413;
      end
      11'b10110000110 : begin
        result = input_1414;
      end
      11'b10110000111 : begin
        result = input_1415;
      end
      11'b10110001000 : begin
        result = input_1416;
      end
      11'b10110001001 : begin
        result = input_1417;
      end
      11'b10110001010 : begin
        result = input_1418;
      end
      11'b10110001011 : begin
        result = input_1419;
      end
      11'b10110001100 : begin
        result = input_1420;
      end
      11'b10110001101 : begin
        result = input_1421;
      end
      11'b10110001110 : begin
        result = input_1422;
      end
      11'b10110001111 : begin
        result = input_1423;
      end
      11'b10110010000 : begin
        result = input_1424;
      end
      11'b10110010001 : begin
        result = input_1425;
      end
      11'b10110010010 : begin
        result = input_1426;
      end
      11'b10110010011 : begin
        result = input_1427;
      end
      11'b10110010100 : begin
        result = input_1428;
      end
      11'b10110010101 : begin
        result = input_1429;
      end
      11'b10110010110 : begin
        result = input_1430;
      end
      11'b10110010111 : begin
        result = input_1431;
      end
      11'b10110011000 : begin
        result = input_1432;
      end
      11'b10110011001 : begin
        result = input_1433;
      end
      11'b10110011010 : begin
        result = input_1434;
      end
      11'b10110011011 : begin
        result = input_1435;
      end
      11'b10110011100 : begin
        result = input_1436;
      end
      11'b10110011101 : begin
        result = input_1437;
      end
      11'b10110011110 : begin
        result = input_1438;
      end
      11'b10110011111 : begin
        result = input_1439;
      end
      11'b10110100000 : begin
        result = input_1440;
      end
      11'b10110100001 : begin
        result = input_1441;
      end
      11'b10110100010 : begin
        result = input_1442;
      end
      11'b10110100011 : begin
        result = input_1443;
      end
      11'b10110100100 : begin
        result = input_1444;
      end
      11'b10110100101 : begin
        result = input_1445;
      end
      11'b10110100110 : begin
        result = input_1446;
      end
      11'b10110100111 : begin
        result = input_1447;
      end
      11'b10110101000 : begin
        result = input_1448;
      end
      11'b10110101001 : begin
        result = input_1449;
      end
      11'b10110101010 : begin
        result = input_1450;
      end
      11'b10110101011 : begin
        result = input_1451;
      end
      11'b10110101100 : begin
        result = input_1452;
      end
      11'b10110101101 : begin
        result = input_1453;
      end
      11'b10110101110 : begin
        result = input_1454;
      end
      11'b10110101111 : begin
        result = input_1455;
      end
      11'b10110110000 : begin
        result = input_1456;
      end
      11'b10110110001 : begin
        result = input_1457;
      end
      11'b10110110010 : begin
        result = input_1458;
      end
      11'b10110110011 : begin
        result = input_1459;
      end
      11'b10110110100 : begin
        result = input_1460;
      end
      11'b10110110101 : begin
        result = input_1461;
      end
      11'b10110110110 : begin
        result = input_1462;
      end
      11'b10110110111 : begin
        result = input_1463;
      end
      11'b10110111000 : begin
        result = input_1464;
      end
      11'b10110111001 : begin
        result = input_1465;
      end
      11'b10110111010 : begin
        result = input_1466;
      end
      11'b10110111011 : begin
        result = input_1467;
      end
      11'b10110111100 : begin
        result = input_1468;
      end
      11'b10110111101 : begin
        result = input_1469;
      end
      11'b10110111110 : begin
        result = input_1470;
      end
      11'b10110111111 : begin
        result = input_1471;
      end
      11'b10111000000 : begin
        result = input_1472;
      end
      11'b10111000001 : begin
        result = input_1473;
      end
      11'b10111000010 : begin
        result = input_1474;
      end
      11'b10111000011 : begin
        result = input_1475;
      end
      11'b10111000100 : begin
        result = input_1476;
      end
      11'b10111000101 : begin
        result = input_1477;
      end
      11'b10111000110 : begin
        result = input_1478;
      end
      11'b10111000111 : begin
        result = input_1479;
      end
      11'b10111001000 : begin
        result = input_1480;
      end
      11'b10111001001 : begin
        result = input_1481;
      end
      11'b10111001010 : begin
        result = input_1482;
      end
      11'b10111001011 : begin
        result = input_1483;
      end
      11'b10111001100 : begin
        result = input_1484;
      end
      11'b10111001101 : begin
        result = input_1485;
      end
      11'b10111001110 : begin
        result = input_1486;
      end
      11'b10111001111 : begin
        result = input_1487;
      end
      11'b10111010000 : begin
        result = input_1488;
      end
      11'b10111010001 : begin
        result = input_1489;
      end
      11'b10111010010 : begin
        result = input_1490;
      end
      11'b10111010011 : begin
        result = input_1491;
      end
      11'b10111010100 : begin
        result = input_1492;
      end
      11'b10111010101 : begin
        result = input_1493;
      end
      11'b10111010110 : begin
        result = input_1494;
      end
      11'b10111010111 : begin
        result = input_1495;
      end
      11'b10111011000 : begin
        result = input_1496;
      end
      11'b10111011001 : begin
        result = input_1497;
      end
      11'b10111011010 : begin
        result = input_1498;
      end
      11'b10111011011 : begin
        result = input_1499;
      end
      11'b10111011100 : begin
        result = input_1500;
      end
      11'b10111011101 : begin
        result = input_1501;
      end
      11'b10111011110 : begin
        result = input_1502;
      end
      11'b10111011111 : begin
        result = input_1503;
      end
      11'b10111100000 : begin
        result = input_1504;
      end
      11'b10111100001 : begin
        result = input_1505;
      end
      11'b10111100010 : begin
        result = input_1506;
      end
      11'b10111100011 : begin
        result = input_1507;
      end
      11'b10111100100 : begin
        result = input_1508;
      end
      11'b10111100101 : begin
        result = input_1509;
      end
      11'b10111100110 : begin
        result = input_1510;
      end
      11'b10111100111 : begin
        result = input_1511;
      end
      11'b10111101000 : begin
        result = input_1512;
      end
      11'b10111101001 : begin
        result = input_1513;
      end
      11'b10111101010 : begin
        result = input_1514;
      end
      11'b10111101011 : begin
        result = input_1515;
      end
      11'b10111101100 : begin
        result = input_1516;
      end
      11'b10111101101 : begin
        result = input_1517;
      end
      11'b10111101110 : begin
        result = input_1518;
      end
      11'b10111101111 : begin
        result = input_1519;
      end
      11'b10111110000 : begin
        result = input_1520;
      end
      11'b10111110001 : begin
        result = input_1521;
      end
      11'b10111110010 : begin
        result = input_1522;
      end
      11'b10111110011 : begin
        result = input_1523;
      end
      11'b10111110100 : begin
        result = input_1524;
      end
      11'b10111110101 : begin
        result = input_1525;
      end
      11'b10111110110 : begin
        result = input_1526;
      end
      11'b10111110111 : begin
        result = input_1527;
      end
      11'b10111111000 : begin
        result = input_1528;
      end
      11'b10111111001 : begin
        result = input_1529;
      end
      11'b10111111010 : begin
        result = input_1530;
      end
      11'b10111111011 : begin
        result = input_1531;
      end
      11'b10111111100 : begin
        result = input_1532;
      end
      11'b10111111101 : begin
        result = input_1533;
      end
      11'b10111111110 : begin
        result = input_1534;
      end
      11'b10111111111 : begin
        result = input_1535;
      end
      11'b11000000000 : begin
        result = input_1536;
      end
      11'b11000000001 : begin
        result = input_1537;
      end
      11'b11000000010 : begin
        result = input_1538;
      end
      11'b11000000011 : begin
        result = input_1539;
      end
      11'b11000000100 : begin
        result = input_1540;
      end
      11'b11000000101 : begin
        result = input_1541;
      end
      11'b11000000110 : begin
        result = input_1542;
      end
      11'b11000000111 : begin
        result = input_1543;
      end
      11'b11000001000 : begin
        result = input_1544;
      end
      11'b11000001001 : begin
        result = input_1545;
      end
      11'b11000001010 : begin
        result = input_1546;
      end
      11'b11000001011 : begin
        result = input_1547;
      end
      11'b11000001100 : begin
        result = input_1548;
      end
      11'b11000001101 : begin
        result = input_1549;
      end
      11'b11000001110 : begin
        result = input_1550;
      end
      11'b11000001111 : begin
        result = input_1551;
      end
      11'b11000010000 : begin
        result = input_1552;
      end
      11'b11000010001 : begin
        result = input_1553;
      end
      11'b11000010010 : begin
        result = input_1554;
      end
      11'b11000010011 : begin
        result = input_1555;
      end
      11'b11000010100 : begin
        result = input_1556;
      end
      11'b11000010101 : begin
        result = input_1557;
      end
      11'b11000010110 : begin
        result = input_1558;
      end
      11'b11000010111 : begin
        result = input_1559;
      end
      11'b11000011000 : begin
        result = input_1560;
      end
      11'b11000011001 : begin
        result = input_1561;
      end
      11'b11000011010 : begin
        result = input_1562;
      end
      11'b11000011011 : begin
        result = input_1563;
      end
      11'b11000011100 : begin
        result = input_1564;
      end
      11'b11000011101 : begin
        result = input_1565;
      end
      11'b11000011110 : begin
        result = input_1566;
      end
      11'b11000011111 : begin
        result = input_1567;
      end
      11'b11000100000 : begin
        result = input_1568;
      end
      11'b11000100001 : begin
        result = input_1569;
      end
      11'b11000100010 : begin
        result = input_1570;
      end
      11'b11000100011 : begin
        result = input_1571;
      end
      11'b11000100100 : begin
        result = input_1572;
      end
      11'b11000100101 : begin
        result = input_1573;
      end
      11'b11000100110 : begin
        result = input_1574;
      end
      11'b11000100111 : begin
        result = input_1575;
      end
      11'b11000101000 : begin
        result = input_1576;
      end
      11'b11000101001 : begin
        result = input_1577;
      end
      11'b11000101010 : begin
        result = input_1578;
      end
      11'b11000101011 : begin
        result = input_1579;
      end
      11'b11000101100 : begin
        result = input_1580;
      end
      11'b11000101101 : begin
        result = input_1581;
      end
      11'b11000101110 : begin
        result = input_1582;
      end
      11'b11000101111 : begin
        result = input_1583;
      end
      11'b11000110000 : begin
        result = input_1584;
      end
      11'b11000110001 : begin
        result = input_1585;
      end
      11'b11000110010 : begin
        result = input_1586;
      end
      11'b11000110011 : begin
        result = input_1587;
      end
      11'b11000110100 : begin
        result = input_1588;
      end
      11'b11000110101 : begin
        result = input_1589;
      end
      11'b11000110110 : begin
        result = input_1590;
      end
      11'b11000110111 : begin
        result = input_1591;
      end
      11'b11000111000 : begin
        result = input_1592;
      end
      11'b11000111001 : begin
        result = input_1593;
      end
      11'b11000111010 : begin
        result = input_1594;
      end
      11'b11000111011 : begin
        result = input_1595;
      end
      11'b11000111100 : begin
        result = input_1596;
      end
      11'b11000111101 : begin
        result = input_1597;
      end
      11'b11000111110 : begin
        result = input_1598;
      end
      11'b11000111111 : begin
        result = input_1599;
      end
      11'b11001000000 : begin
        result = input_1600;
      end
      11'b11001000001 : begin
        result = input_1601;
      end
      11'b11001000010 : begin
        result = input_1602;
      end
      11'b11001000011 : begin
        result = input_1603;
      end
      11'b11001000100 : begin
        result = input_1604;
      end
      11'b11001000101 : begin
        result = input_1605;
      end
      11'b11001000110 : begin
        result = input_1606;
      end
      11'b11001000111 : begin
        result = input_1607;
      end
      11'b11001001000 : begin
        result = input_1608;
      end
      11'b11001001001 : begin
        result = input_1609;
      end
      11'b11001001010 : begin
        result = input_1610;
      end
      11'b11001001011 : begin
        result = input_1611;
      end
      11'b11001001100 : begin
        result = input_1612;
      end
      11'b11001001101 : begin
        result = input_1613;
      end
      11'b11001001110 : begin
        result = input_1614;
      end
      11'b11001001111 : begin
        result = input_1615;
      end
      11'b11001010000 : begin
        result = input_1616;
      end
      11'b11001010001 : begin
        result = input_1617;
      end
      11'b11001010010 : begin
        result = input_1618;
      end
      11'b11001010011 : begin
        result = input_1619;
      end
      11'b11001010100 : begin
        result = input_1620;
      end
      11'b11001010101 : begin
        result = input_1621;
      end
      11'b11001010110 : begin
        result = input_1622;
      end
      11'b11001010111 : begin
        result = input_1623;
      end
      11'b11001011000 : begin
        result = input_1624;
      end
      11'b11001011001 : begin
        result = input_1625;
      end
      11'b11001011010 : begin
        result = input_1626;
      end
      11'b11001011011 : begin
        result = input_1627;
      end
      11'b11001011100 : begin
        result = input_1628;
      end
      11'b11001011101 : begin
        result = input_1629;
      end
      11'b11001011110 : begin
        result = input_1630;
      end
      11'b11001011111 : begin
        result = input_1631;
      end
      11'b11001100000 : begin
        result = input_1632;
      end
      11'b11001100001 : begin
        result = input_1633;
      end
      11'b11001100010 : begin
        result = input_1634;
      end
      11'b11001100011 : begin
        result = input_1635;
      end
      11'b11001100100 : begin
        result = input_1636;
      end
      11'b11001100101 : begin
        result = input_1637;
      end
      11'b11001100110 : begin
        result = input_1638;
      end
      11'b11001100111 : begin
        result = input_1639;
      end
      11'b11001101000 : begin
        result = input_1640;
      end
      11'b11001101001 : begin
        result = input_1641;
      end
      11'b11001101010 : begin
        result = input_1642;
      end
      11'b11001101011 : begin
        result = input_1643;
      end
      11'b11001101100 : begin
        result = input_1644;
      end
      11'b11001101101 : begin
        result = input_1645;
      end
      11'b11001101110 : begin
        result = input_1646;
      end
      11'b11001101111 : begin
        result = input_1647;
      end
      11'b11001110000 : begin
        result = input_1648;
      end
      11'b11001110001 : begin
        result = input_1649;
      end
      11'b11001110010 : begin
        result = input_1650;
      end
      11'b11001110011 : begin
        result = input_1651;
      end
      11'b11001110100 : begin
        result = input_1652;
      end
      11'b11001110101 : begin
        result = input_1653;
      end
      11'b11001110110 : begin
        result = input_1654;
      end
      11'b11001110111 : begin
        result = input_1655;
      end
      11'b11001111000 : begin
        result = input_1656;
      end
      11'b11001111001 : begin
        result = input_1657;
      end
      11'b11001111010 : begin
        result = input_1658;
      end
      11'b11001111011 : begin
        result = input_1659;
      end
      11'b11001111100 : begin
        result = input_1660;
      end
      11'b11001111101 : begin
        result = input_1661;
      end
      11'b11001111110 : begin
        result = input_1662;
      end
      11'b11001111111 : begin
        result = input_1663;
      end
      11'b11010000000 : begin
        result = input_1664;
      end
      11'b11010000001 : begin
        result = input_1665;
      end
      11'b11010000010 : begin
        result = input_1666;
      end
      11'b11010000011 : begin
        result = input_1667;
      end
      11'b11010000100 : begin
        result = input_1668;
      end
      11'b11010000101 : begin
        result = input_1669;
      end
      11'b11010000110 : begin
        result = input_1670;
      end
      11'b11010000111 : begin
        result = input_1671;
      end
      11'b11010001000 : begin
        result = input_1672;
      end
      11'b11010001001 : begin
        result = input_1673;
      end
      11'b11010001010 : begin
        result = input_1674;
      end
      11'b11010001011 : begin
        result = input_1675;
      end
      11'b11010001100 : begin
        result = input_1676;
      end
      11'b11010001101 : begin
        result = input_1677;
      end
      11'b11010001110 : begin
        result = input_1678;
      end
      11'b11010001111 : begin
        result = input_1679;
      end
      11'b11010010000 : begin
        result = input_1680;
      end
      11'b11010010001 : begin
        result = input_1681;
      end
      11'b11010010010 : begin
        result = input_1682;
      end
      11'b11010010011 : begin
        result = input_1683;
      end
      11'b11010010100 : begin
        result = input_1684;
      end
      11'b11010010101 : begin
        result = input_1685;
      end
      11'b11010010110 : begin
        result = input_1686;
      end
      11'b11010010111 : begin
        result = input_1687;
      end
      11'b11010011000 : begin
        result = input_1688;
      end
      11'b11010011001 : begin
        result = input_1689;
      end
      11'b11010011010 : begin
        result = input_1690;
      end
      11'b11010011011 : begin
        result = input_1691;
      end
      11'b11010011100 : begin
        result = input_1692;
      end
      11'b11010011101 : begin
        result = input_1693;
      end
      11'b11010011110 : begin
        result = input_1694;
      end
      11'b11010011111 : begin
        result = input_1695;
      end
      11'b11010100000 : begin
        result = input_1696;
      end
      11'b11010100001 : begin
        result = input_1697;
      end
      11'b11010100010 : begin
        result = input_1698;
      end
      11'b11010100011 : begin
        result = input_1699;
      end
      11'b11010100100 : begin
        result = input_1700;
      end
      11'b11010100101 : begin
        result = input_1701;
      end
      11'b11010100110 : begin
        result = input_1702;
      end
      11'b11010100111 : begin
        result = input_1703;
      end
      11'b11010101000 : begin
        result = input_1704;
      end
      11'b11010101001 : begin
        result = input_1705;
      end
      11'b11010101010 : begin
        result = input_1706;
      end
      11'b11010101011 : begin
        result = input_1707;
      end
      11'b11010101100 : begin
        result = input_1708;
      end
      11'b11010101101 : begin
        result = input_1709;
      end
      11'b11010101110 : begin
        result = input_1710;
      end
      11'b11010101111 : begin
        result = input_1711;
      end
      11'b11010110000 : begin
        result = input_1712;
      end
      11'b11010110001 : begin
        result = input_1713;
      end
      11'b11010110010 : begin
        result = input_1714;
      end
      11'b11010110011 : begin
        result = input_1715;
      end
      11'b11010110100 : begin
        result = input_1716;
      end
      11'b11010110101 : begin
        result = input_1717;
      end
      11'b11010110110 : begin
        result = input_1718;
      end
      11'b11010110111 : begin
        result = input_1719;
      end
      11'b11010111000 : begin
        result = input_1720;
      end
      11'b11010111001 : begin
        result = input_1721;
      end
      11'b11010111010 : begin
        result = input_1722;
      end
      11'b11010111011 : begin
        result = input_1723;
      end
      11'b11010111100 : begin
        result = input_1724;
      end
      11'b11010111101 : begin
        result = input_1725;
      end
      11'b11010111110 : begin
        result = input_1726;
      end
      11'b11010111111 : begin
        result = input_1727;
      end
      11'b11011000000 : begin
        result = input_1728;
      end
      11'b11011000001 : begin
        result = input_1729;
      end
      11'b11011000010 : begin
        result = input_1730;
      end
      11'b11011000011 : begin
        result = input_1731;
      end
      11'b11011000100 : begin
        result = input_1732;
      end
      11'b11011000101 : begin
        result = input_1733;
      end
      11'b11011000110 : begin
        result = input_1734;
      end
      11'b11011000111 : begin
        result = input_1735;
      end
      11'b11011001000 : begin
        result = input_1736;
      end
      11'b11011001001 : begin
        result = input_1737;
      end
      11'b11011001010 : begin
        result = input_1738;
      end
      11'b11011001011 : begin
        result = input_1739;
      end
      11'b11011001100 : begin
        result = input_1740;
      end
      11'b11011001101 : begin
        result = input_1741;
      end
      11'b11011001110 : begin
        result = input_1742;
      end
      11'b11011001111 : begin
        result = input_1743;
      end
      11'b11011010000 : begin
        result = input_1744;
      end
      11'b11011010001 : begin
        result = input_1745;
      end
      11'b11011010010 : begin
        result = input_1746;
      end
      11'b11011010011 : begin
        result = input_1747;
      end
      11'b11011010100 : begin
        result = input_1748;
      end
      11'b11011010101 : begin
        result = input_1749;
      end
      11'b11011010110 : begin
        result = input_1750;
      end
      11'b11011010111 : begin
        result = input_1751;
      end
      11'b11011011000 : begin
        result = input_1752;
      end
      11'b11011011001 : begin
        result = input_1753;
      end
      11'b11011011010 : begin
        result = input_1754;
      end
      11'b11011011011 : begin
        result = input_1755;
      end
      11'b11011011100 : begin
        result = input_1756;
      end
      11'b11011011101 : begin
        result = input_1757;
      end
      11'b11011011110 : begin
        result = input_1758;
      end
      11'b11011011111 : begin
        result = input_1759;
      end
      11'b11011100000 : begin
        result = input_1760;
      end
      11'b11011100001 : begin
        result = input_1761;
      end
      11'b11011100010 : begin
        result = input_1762;
      end
      11'b11011100011 : begin
        result = input_1763;
      end
      11'b11011100100 : begin
        result = input_1764;
      end
      11'b11011100101 : begin
        result = input_1765;
      end
      11'b11011100110 : begin
        result = input_1766;
      end
      11'b11011100111 : begin
        result = input_1767;
      end
      11'b11011101000 : begin
        result = input_1768;
      end
      11'b11011101001 : begin
        result = input_1769;
      end
      11'b11011101010 : begin
        result = input_1770;
      end
      11'b11011101011 : begin
        result = input_1771;
      end
      11'b11011101100 : begin
        result = input_1772;
      end
      11'b11011101101 : begin
        result = input_1773;
      end
      11'b11011101110 : begin
        result = input_1774;
      end
      11'b11011101111 : begin
        result = input_1775;
      end
      11'b11011110000 : begin
        result = input_1776;
      end
      11'b11011110001 : begin
        result = input_1777;
      end
      11'b11011110010 : begin
        result = input_1778;
      end
      11'b11011110011 : begin
        result = input_1779;
      end
      11'b11011110100 : begin
        result = input_1780;
      end
      11'b11011110101 : begin
        result = input_1781;
      end
      11'b11011110110 : begin
        result = input_1782;
      end
      11'b11011110111 : begin
        result = input_1783;
      end
      11'b11011111000 : begin
        result = input_1784;
      end
      11'b11011111001 : begin
        result = input_1785;
      end
      11'b11011111010 : begin
        result = input_1786;
      end
      11'b11011111011 : begin
        result = input_1787;
      end
      11'b11011111100 : begin
        result = input_1788;
      end
      11'b11011111101 : begin
        result = input_1789;
      end
      11'b11011111110 : begin
        result = input_1790;
      end
      default : begin
        result = input_1791;
      end
    endcase
    MUX_v_16_1792_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_384_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [15:0] input_56;
    input [15:0] input_57;
    input [15:0] input_58;
    input [15:0] input_59;
    input [15:0] input_60;
    input [15:0] input_61;
    input [15:0] input_62;
    input [15:0] input_63;
    input [15:0] input_64;
    input [15:0] input_65;
    input [15:0] input_66;
    input [15:0] input_67;
    input [15:0] input_68;
    input [15:0] input_69;
    input [15:0] input_70;
    input [15:0] input_71;
    input [15:0] input_72;
    input [15:0] input_73;
    input [15:0] input_74;
    input [15:0] input_75;
    input [15:0] input_76;
    input [15:0] input_77;
    input [15:0] input_78;
    input [15:0] input_79;
    input [15:0] input_80;
    input [15:0] input_81;
    input [15:0] input_82;
    input [15:0] input_83;
    input [15:0] input_84;
    input [15:0] input_85;
    input [15:0] input_86;
    input [15:0] input_87;
    input [15:0] input_88;
    input [15:0] input_89;
    input [15:0] input_90;
    input [15:0] input_91;
    input [15:0] input_92;
    input [15:0] input_93;
    input [15:0] input_94;
    input [15:0] input_95;
    input [15:0] input_96;
    input [15:0] input_97;
    input [15:0] input_98;
    input [15:0] input_99;
    input [15:0] input_100;
    input [15:0] input_101;
    input [15:0] input_102;
    input [15:0] input_103;
    input [15:0] input_104;
    input [15:0] input_105;
    input [15:0] input_106;
    input [15:0] input_107;
    input [15:0] input_108;
    input [15:0] input_109;
    input [15:0] input_110;
    input [15:0] input_111;
    input [15:0] input_112;
    input [15:0] input_113;
    input [15:0] input_114;
    input [15:0] input_115;
    input [15:0] input_116;
    input [15:0] input_117;
    input [15:0] input_118;
    input [15:0] input_119;
    input [15:0] input_120;
    input [15:0] input_121;
    input [15:0] input_122;
    input [15:0] input_123;
    input [15:0] input_124;
    input [15:0] input_125;
    input [15:0] input_126;
    input [15:0] input_127;
    input [15:0] input_128;
    input [15:0] input_129;
    input [15:0] input_130;
    input [15:0] input_131;
    input [15:0] input_132;
    input [15:0] input_133;
    input [15:0] input_134;
    input [15:0] input_135;
    input [15:0] input_136;
    input [15:0] input_137;
    input [15:0] input_138;
    input [15:0] input_139;
    input [15:0] input_140;
    input [15:0] input_141;
    input [15:0] input_142;
    input [15:0] input_143;
    input [15:0] input_144;
    input [15:0] input_145;
    input [15:0] input_146;
    input [15:0] input_147;
    input [15:0] input_148;
    input [15:0] input_149;
    input [15:0] input_150;
    input [15:0] input_151;
    input [15:0] input_152;
    input [15:0] input_153;
    input [15:0] input_154;
    input [15:0] input_155;
    input [15:0] input_156;
    input [15:0] input_157;
    input [15:0] input_158;
    input [15:0] input_159;
    input [15:0] input_160;
    input [15:0] input_161;
    input [15:0] input_162;
    input [15:0] input_163;
    input [15:0] input_164;
    input [15:0] input_165;
    input [15:0] input_166;
    input [15:0] input_167;
    input [15:0] input_168;
    input [15:0] input_169;
    input [15:0] input_170;
    input [15:0] input_171;
    input [15:0] input_172;
    input [15:0] input_173;
    input [15:0] input_174;
    input [15:0] input_175;
    input [15:0] input_176;
    input [15:0] input_177;
    input [15:0] input_178;
    input [15:0] input_179;
    input [15:0] input_180;
    input [15:0] input_181;
    input [15:0] input_182;
    input [15:0] input_183;
    input [15:0] input_184;
    input [15:0] input_185;
    input [15:0] input_186;
    input [15:0] input_187;
    input [15:0] input_188;
    input [15:0] input_189;
    input [15:0] input_190;
    input [15:0] input_191;
    input [15:0] input_192;
    input [15:0] input_193;
    input [15:0] input_194;
    input [15:0] input_195;
    input [15:0] input_196;
    input [15:0] input_197;
    input [15:0] input_198;
    input [15:0] input_199;
    input [15:0] input_200;
    input [15:0] input_201;
    input [15:0] input_202;
    input [15:0] input_203;
    input [15:0] input_204;
    input [15:0] input_205;
    input [15:0] input_206;
    input [15:0] input_207;
    input [15:0] input_208;
    input [15:0] input_209;
    input [15:0] input_210;
    input [15:0] input_211;
    input [15:0] input_212;
    input [15:0] input_213;
    input [15:0] input_214;
    input [15:0] input_215;
    input [15:0] input_216;
    input [15:0] input_217;
    input [15:0] input_218;
    input [15:0] input_219;
    input [15:0] input_220;
    input [15:0] input_221;
    input [15:0] input_222;
    input [15:0] input_223;
    input [15:0] input_224;
    input [15:0] input_225;
    input [15:0] input_226;
    input [15:0] input_227;
    input [15:0] input_228;
    input [15:0] input_229;
    input [15:0] input_230;
    input [15:0] input_231;
    input [15:0] input_232;
    input [15:0] input_233;
    input [15:0] input_234;
    input [15:0] input_235;
    input [15:0] input_236;
    input [15:0] input_237;
    input [15:0] input_238;
    input [15:0] input_239;
    input [15:0] input_240;
    input [15:0] input_241;
    input [15:0] input_242;
    input [15:0] input_243;
    input [15:0] input_244;
    input [15:0] input_245;
    input [15:0] input_246;
    input [15:0] input_247;
    input [15:0] input_248;
    input [15:0] input_249;
    input [15:0] input_250;
    input [15:0] input_251;
    input [15:0] input_252;
    input [15:0] input_253;
    input [15:0] input_254;
    input [15:0] input_255;
    input [15:0] input_256;
    input [15:0] input_257;
    input [15:0] input_258;
    input [15:0] input_259;
    input [15:0] input_260;
    input [15:0] input_261;
    input [15:0] input_262;
    input [15:0] input_263;
    input [15:0] input_264;
    input [15:0] input_265;
    input [15:0] input_266;
    input [15:0] input_267;
    input [15:0] input_268;
    input [15:0] input_269;
    input [15:0] input_270;
    input [15:0] input_271;
    input [15:0] input_272;
    input [15:0] input_273;
    input [15:0] input_274;
    input [15:0] input_275;
    input [15:0] input_276;
    input [15:0] input_277;
    input [15:0] input_278;
    input [15:0] input_279;
    input [15:0] input_280;
    input [15:0] input_281;
    input [15:0] input_282;
    input [15:0] input_283;
    input [15:0] input_284;
    input [15:0] input_285;
    input [15:0] input_286;
    input [15:0] input_287;
    input [15:0] input_288;
    input [15:0] input_289;
    input [15:0] input_290;
    input [15:0] input_291;
    input [15:0] input_292;
    input [15:0] input_293;
    input [15:0] input_294;
    input [15:0] input_295;
    input [15:0] input_296;
    input [15:0] input_297;
    input [15:0] input_298;
    input [15:0] input_299;
    input [15:0] input_300;
    input [15:0] input_301;
    input [15:0] input_302;
    input [15:0] input_303;
    input [15:0] input_304;
    input [15:0] input_305;
    input [15:0] input_306;
    input [15:0] input_307;
    input [15:0] input_308;
    input [15:0] input_309;
    input [15:0] input_310;
    input [15:0] input_311;
    input [15:0] input_312;
    input [15:0] input_313;
    input [15:0] input_314;
    input [15:0] input_315;
    input [15:0] input_316;
    input [15:0] input_317;
    input [15:0] input_318;
    input [15:0] input_319;
    input [15:0] input_320;
    input [15:0] input_321;
    input [15:0] input_322;
    input [15:0] input_323;
    input [15:0] input_324;
    input [15:0] input_325;
    input [15:0] input_326;
    input [15:0] input_327;
    input [15:0] input_328;
    input [15:0] input_329;
    input [15:0] input_330;
    input [15:0] input_331;
    input [15:0] input_332;
    input [15:0] input_333;
    input [15:0] input_334;
    input [15:0] input_335;
    input [15:0] input_336;
    input [15:0] input_337;
    input [15:0] input_338;
    input [15:0] input_339;
    input [15:0] input_340;
    input [15:0] input_341;
    input [15:0] input_342;
    input [15:0] input_343;
    input [15:0] input_344;
    input [15:0] input_345;
    input [15:0] input_346;
    input [15:0] input_347;
    input [15:0] input_348;
    input [15:0] input_349;
    input [15:0] input_350;
    input [15:0] input_351;
    input [15:0] input_352;
    input [15:0] input_353;
    input [15:0] input_354;
    input [15:0] input_355;
    input [15:0] input_356;
    input [15:0] input_357;
    input [15:0] input_358;
    input [15:0] input_359;
    input [15:0] input_360;
    input [15:0] input_361;
    input [15:0] input_362;
    input [15:0] input_363;
    input [15:0] input_364;
    input [15:0] input_365;
    input [15:0] input_366;
    input [15:0] input_367;
    input [15:0] input_368;
    input [15:0] input_369;
    input [15:0] input_370;
    input [15:0] input_371;
    input [15:0] input_372;
    input [15:0] input_373;
    input [15:0] input_374;
    input [15:0] input_375;
    input [15:0] input_376;
    input [15:0] input_377;
    input [15:0] input_378;
    input [15:0] input_379;
    input [15:0] input_380;
    input [15:0] input_381;
    input [15:0] input_382;
    input [15:0] input_383;
    input [8:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = input_0;
      end
      9'b000000001 : begin
        result = input_1;
      end
      9'b000000010 : begin
        result = input_2;
      end
      9'b000000011 : begin
        result = input_3;
      end
      9'b000000100 : begin
        result = input_4;
      end
      9'b000000101 : begin
        result = input_5;
      end
      9'b000000110 : begin
        result = input_6;
      end
      9'b000000111 : begin
        result = input_7;
      end
      9'b000001000 : begin
        result = input_8;
      end
      9'b000001001 : begin
        result = input_9;
      end
      9'b000001010 : begin
        result = input_10;
      end
      9'b000001011 : begin
        result = input_11;
      end
      9'b000001100 : begin
        result = input_12;
      end
      9'b000001101 : begin
        result = input_13;
      end
      9'b000001110 : begin
        result = input_14;
      end
      9'b000001111 : begin
        result = input_15;
      end
      9'b000010000 : begin
        result = input_16;
      end
      9'b000010001 : begin
        result = input_17;
      end
      9'b000010010 : begin
        result = input_18;
      end
      9'b000010011 : begin
        result = input_19;
      end
      9'b000010100 : begin
        result = input_20;
      end
      9'b000010101 : begin
        result = input_21;
      end
      9'b000010110 : begin
        result = input_22;
      end
      9'b000010111 : begin
        result = input_23;
      end
      9'b000011000 : begin
        result = input_24;
      end
      9'b000011001 : begin
        result = input_25;
      end
      9'b000011010 : begin
        result = input_26;
      end
      9'b000011011 : begin
        result = input_27;
      end
      9'b000011100 : begin
        result = input_28;
      end
      9'b000011101 : begin
        result = input_29;
      end
      9'b000011110 : begin
        result = input_30;
      end
      9'b000011111 : begin
        result = input_31;
      end
      9'b000100000 : begin
        result = input_32;
      end
      9'b000100001 : begin
        result = input_33;
      end
      9'b000100010 : begin
        result = input_34;
      end
      9'b000100011 : begin
        result = input_35;
      end
      9'b000100100 : begin
        result = input_36;
      end
      9'b000100101 : begin
        result = input_37;
      end
      9'b000100110 : begin
        result = input_38;
      end
      9'b000100111 : begin
        result = input_39;
      end
      9'b000101000 : begin
        result = input_40;
      end
      9'b000101001 : begin
        result = input_41;
      end
      9'b000101010 : begin
        result = input_42;
      end
      9'b000101011 : begin
        result = input_43;
      end
      9'b000101100 : begin
        result = input_44;
      end
      9'b000101101 : begin
        result = input_45;
      end
      9'b000101110 : begin
        result = input_46;
      end
      9'b000101111 : begin
        result = input_47;
      end
      9'b000110000 : begin
        result = input_48;
      end
      9'b000110001 : begin
        result = input_49;
      end
      9'b000110010 : begin
        result = input_50;
      end
      9'b000110011 : begin
        result = input_51;
      end
      9'b000110100 : begin
        result = input_52;
      end
      9'b000110101 : begin
        result = input_53;
      end
      9'b000110110 : begin
        result = input_54;
      end
      9'b000110111 : begin
        result = input_55;
      end
      9'b000111000 : begin
        result = input_56;
      end
      9'b000111001 : begin
        result = input_57;
      end
      9'b000111010 : begin
        result = input_58;
      end
      9'b000111011 : begin
        result = input_59;
      end
      9'b000111100 : begin
        result = input_60;
      end
      9'b000111101 : begin
        result = input_61;
      end
      9'b000111110 : begin
        result = input_62;
      end
      9'b000111111 : begin
        result = input_63;
      end
      9'b001000000 : begin
        result = input_64;
      end
      9'b001000001 : begin
        result = input_65;
      end
      9'b001000010 : begin
        result = input_66;
      end
      9'b001000011 : begin
        result = input_67;
      end
      9'b001000100 : begin
        result = input_68;
      end
      9'b001000101 : begin
        result = input_69;
      end
      9'b001000110 : begin
        result = input_70;
      end
      9'b001000111 : begin
        result = input_71;
      end
      9'b001001000 : begin
        result = input_72;
      end
      9'b001001001 : begin
        result = input_73;
      end
      9'b001001010 : begin
        result = input_74;
      end
      9'b001001011 : begin
        result = input_75;
      end
      9'b001001100 : begin
        result = input_76;
      end
      9'b001001101 : begin
        result = input_77;
      end
      9'b001001110 : begin
        result = input_78;
      end
      9'b001001111 : begin
        result = input_79;
      end
      9'b001010000 : begin
        result = input_80;
      end
      9'b001010001 : begin
        result = input_81;
      end
      9'b001010010 : begin
        result = input_82;
      end
      9'b001010011 : begin
        result = input_83;
      end
      9'b001010100 : begin
        result = input_84;
      end
      9'b001010101 : begin
        result = input_85;
      end
      9'b001010110 : begin
        result = input_86;
      end
      9'b001010111 : begin
        result = input_87;
      end
      9'b001011000 : begin
        result = input_88;
      end
      9'b001011001 : begin
        result = input_89;
      end
      9'b001011010 : begin
        result = input_90;
      end
      9'b001011011 : begin
        result = input_91;
      end
      9'b001011100 : begin
        result = input_92;
      end
      9'b001011101 : begin
        result = input_93;
      end
      9'b001011110 : begin
        result = input_94;
      end
      9'b001011111 : begin
        result = input_95;
      end
      9'b001100000 : begin
        result = input_96;
      end
      9'b001100001 : begin
        result = input_97;
      end
      9'b001100010 : begin
        result = input_98;
      end
      9'b001100011 : begin
        result = input_99;
      end
      9'b001100100 : begin
        result = input_100;
      end
      9'b001100101 : begin
        result = input_101;
      end
      9'b001100110 : begin
        result = input_102;
      end
      9'b001100111 : begin
        result = input_103;
      end
      9'b001101000 : begin
        result = input_104;
      end
      9'b001101001 : begin
        result = input_105;
      end
      9'b001101010 : begin
        result = input_106;
      end
      9'b001101011 : begin
        result = input_107;
      end
      9'b001101100 : begin
        result = input_108;
      end
      9'b001101101 : begin
        result = input_109;
      end
      9'b001101110 : begin
        result = input_110;
      end
      9'b001101111 : begin
        result = input_111;
      end
      9'b001110000 : begin
        result = input_112;
      end
      9'b001110001 : begin
        result = input_113;
      end
      9'b001110010 : begin
        result = input_114;
      end
      9'b001110011 : begin
        result = input_115;
      end
      9'b001110100 : begin
        result = input_116;
      end
      9'b001110101 : begin
        result = input_117;
      end
      9'b001110110 : begin
        result = input_118;
      end
      9'b001110111 : begin
        result = input_119;
      end
      9'b001111000 : begin
        result = input_120;
      end
      9'b001111001 : begin
        result = input_121;
      end
      9'b001111010 : begin
        result = input_122;
      end
      9'b001111011 : begin
        result = input_123;
      end
      9'b001111100 : begin
        result = input_124;
      end
      9'b001111101 : begin
        result = input_125;
      end
      9'b001111110 : begin
        result = input_126;
      end
      9'b001111111 : begin
        result = input_127;
      end
      9'b010000000 : begin
        result = input_128;
      end
      9'b010000001 : begin
        result = input_129;
      end
      9'b010000010 : begin
        result = input_130;
      end
      9'b010000011 : begin
        result = input_131;
      end
      9'b010000100 : begin
        result = input_132;
      end
      9'b010000101 : begin
        result = input_133;
      end
      9'b010000110 : begin
        result = input_134;
      end
      9'b010000111 : begin
        result = input_135;
      end
      9'b010001000 : begin
        result = input_136;
      end
      9'b010001001 : begin
        result = input_137;
      end
      9'b010001010 : begin
        result = input_138;
      end
      9'b010001011 : begin
        result = input_139;
      end
      9'b010001100 : begin
        result = input_140;
      end
      9'b010001101 : begin
        result = input_141;
      end
      9'b010001110 : begin
        result = input_142;
      end
      9'b010001111 : begin
        result = input_143;
      end
      9'b010010000 : begin
        result = input_144;
      end
      9'b010010001 : begin
        result = input_145;
      end
      9'b010010010 : begin
        result = input_146;
      end
      9'b010010011 : begin
        result = input_147;
      end
      9'b010010100 : begin
        result = input_148;
      end
      9'b010010101 : begin
        result = input_149;
      end
      9'b010010110 : begin
        result = input_150;
      end
      9'b010010111 : begin
        result = input_151;
      end
      9'b010011000 : begin
        result = input_152;
      end
      9'b010011001 : begin
        result = input_153;
      end
      9'b010011010 : begin
        result = input_154;
      end
      9'b010011011 : begin
        result = input_155;
      end
      9'b010011100 : begin
        result = input_156;
      end
      9'b010011101 : begin
        result = input_157;
      end
      9'b010011110 : begin
        result = input_158;
      end
      9'b010011111 : begin
        result = input_159;
      end
      9'b010100000 : begin
        result = input_160;
      end
      9'b010100001 : begin
        result = input_161;
      end
      9'b010100010 : begin
        result = input_162;
      end
      9'b010100011 : begin
        result = input_163;
      end
      9'b010100100 : begin
        result = input_164;
      end
      9'b010100101 : begin
        result = input_165;
      end
      9'b010100110 : begin
        result = input_166;
      end
      9'b010100111 : begin
        result = input_167;
      end
      9'b010101000 : begin
        result = input_168;
      end
      9'b010101001 : begin
        result = input_169;
      end
      9'b010101010 : begin
        result = input_170;
      end
      9'b010101011 : begin
        result = input_171;
      end
      9'b010101100 : begin
        result = input_172;
      end
      9'b010101101 : begin
        result = input_173;
      end
      9'b010101110 : begin
        result = input_174;
      end
      9'b010101111 : begin
        result = input_175;
      end
      9'b010110000 : begin
        result = input_176;
      end
      9'b010110001 : begin
        result = input_177;
      end
      9'b010110010 : begin
        result = input_178;
      end
      9'b010110011 : begin
        result = input_179;
      end
      9'b010110100 : begin
        result = input_180;
      end
      9'b010110101 : begin
        result = input_181;
      end
      9'b010110110 : begin
        result = input_182;
      end
      9'b010110111 : begin
        result = input_183;
      end
      9'b010111000 : begin
        result = input_184;
      end
      9'b010111001 : begin
        result = input_185;
      end
      9'b010111010 : begin
        result = input_186;
      end
      9'b010111011 : begin
        result = input_187;
      end
      9'b010111100 : begin
        result = input_188;
      end
      9'b010111101 : begin
        result = input_189;
      end
      9'b010111110 : begin
        result = input_190;
      end
      9'b010111111 : begin
        result = input_191;
      end
      9'b011000000 : begin
        result = input_192;
      end
      9'b011000001 : begin
        result = input_193;
      end
      9'b011000010 : begin
        result = input_194;
      end
      9'b011000011 : begin
        result = input_195;
      end
      9'b011000100 : begin
        result = input_196;
      end
      9'b011000101 : begin
        result = input_197;
      end
      9'b011000110 : begin
        result = input_198;
      end
      9'b011000111 : begin
        result = input_199;
      end
      9'b011001000 : begin
        result = input_200;
      end
      9'b011001001 : begin
        result = input_201;
      end
      9'b011001010 : begin
        result = input_202;
      end
      9'b011001011 : begin
        result = input_203;
      end
      9'b011001100 : begin
        result = input_204;
      end
      9'b011001101 : begin
        result = input_205;
      end
      9'b011001110 : begin
        result = input_206;
      end
      9'b011001111 : begin
        result = input_207;
      end
      9'b011010000 : begin
        result = input_208;
      end
      9'b011010001 : begin
        result = input_209;
      end
      9'b011010010 : begin
        result = input_210;
      end
      9'b011010011 : begin
        result = input_211;
      end
      9'b011010100 : begin
        result = input_212;
      end
      9'b011010101 : begin
        result = input_213;
      end
      9'b011010110 : begin
        result = input_214;
      end
      9'b011010111 : begin
        result = input_215;
      end
      9'b011011000 : begin
        result = input_216;
      end
      9'b011011001 : begin
        result = input_217;
      end
      9'b011011010 : begin
        result = input_218;
      end
      9'b011011011 : begin
        result = input_219;
      end
      9'b011011100 : begin
        result = input_220;
      end
      9'b011011101 : begin
        result = input_221;
      end
      9'b011011110 : begin
        result = input_222;
      end
      9'b011011111 : begin
        result = input_223;
      end
      9'b011100000 : begin
        result = input_224;
      end
      9'b011100001 : begin
        result = input_225;
      end
      9'b011100010 : begin
        result = input_226;
      end
      9'b011100011 : begin
        result = input_227;
      end
      9'b011100100 : begin
        result = input_228;
      end
      9'b011100101 : begin
        result = input_229;
      end
      9'b011100110 : begin
        result = input_230;
      end
      9'b011100111 : begin
        result = input_231;
      end
      9'b011101000 : begin
        result = input_232;
      end
      9'b011101001 : begin
        result = input_233;
      end
      9'b011101010 : begin
        result = input_234;
      end
      9'b011101011 : begin
        result = input_235;
      end
      9'b011101100 : begin
        result = input_236;
      end
      9'b011101101 : begin
        result = input_237;
      end
      9'b011101110 : begin
        result = input_238;
      end
      9'b011101111 : begin
        result = input_239;
      end
      9'b011110000 : begin
        result = input_240;
      end
      9'b011110001 : begin
        result = input_241;
      end
      9'b011110010 : begin
        result = input_242;
      end
      9'b011110011 : begin
        result = input_243;
      end
      9'b011110100 : begin
        result = input_244;
      end
      9'b011110101 : begin
        result = input_245;
      end
      9'b011110110 : begin
        result = input_246;
      end
      9'b011110111 : begin
        result = input_247;
      end
      9'b011111000 : begin
        result = input_248;
      end
      9'b011111001 : begin
        result = input_249;
      end
      9'b011111010 : begin
        result = input_250;
      end
      9'b011111011 : begin
        result = input_251;
      end
      9'b011111100 : begin
        result = input_252;
      end
      9'b011111101 : begin
        result = input_253;
      end
      9'b011111110 : begin
        result = input_254;
      end
      9'b011111111 : begin
        result = input_255;
      end
      9'b100000000 : begin
        result = input_256;
      end
      9'b100000001 : begin
        result = input_257;
      end
      9'b100000010 : begin
        result = input_258;
      end
      9'b100000011 : begin
        result = input_259;
      end
      9'b100000100 : begin
        result = input_260;
      end
      9'b100000101 : begin
        result = input_261;
      end
      9'b100000110 : begin
        result = input_262;
      end
      9'b100000111 : begin
        result = input_263;
      end
      9'b100001000 : begin
        result = input_264;
      end
      9'b100001001 : begin
        result = input_265;
      end
      9'b100001010 : begin
        result = input_266;
      end
      9'b100001011 : begin
        result = input_267;
      end
      9'b100001100 : begin
        result = input_268;
      end
      9'b100001101 : begin
        result = input_269;
      end
      9'b100001110 : begin
        result = input_270;
      end
      9'b100001111 : begin
        result = input_271;
      end
      9'b100010000 : begin
        result = input_272;
      end
      9'b100010001 : begin
        result = input_273;
      end
      9'b100010010 : begin
        result = input_274;
      end
      9'b100010011 : begin
        result = input_275;
      end
      9'b100010100 : begin
        result = input_276;
      end
      9'b100010101 : begin
        result = input_277;
      end
      9'b100010110 : begin
        result = input_278;
      end
      9'b100010111 : begin
        result = input_279;
      end
      9'b100011000 : begin
        result = input_280;
      end
      9'b100011001 : begin
        result = input_281;
      end
      9'b100011010 : begin
        result = input_282;
      end
      9'b100011011 : begin
        result = input_283;
      end
      9'b100011100 : begin
        result = input_284;
      end
      9'b100011101 : begin
        result = input_285;
      end
      9'b100011110 : begin
        result = input_286;
      end
      9'b100011111 : begin
        result = input_287;
      end
      9'b100100000 : begin
        result = input_288;
      end
      9'b100100001 : begin
        result = input_289;
      end
      9'b100100010 : begin
        result = input_290;
      end
      9'b100100011 : begin
        result = input_291;
      end
      9'b100100100 : begin
        result = input_292;
      end
      9'b100100101 : begin
        result = input_293;
      end
      9'b100100110 : begin
        result = input_294;
      end
      9'b100100111 : begin
        result = input_295;
      end
      9'b100101000 : begin
        result = input_296;
      end
      9'b100101001 : begin
        result = input_297;
      end
      9'b100101010 : begin
        result = input_298;
      end
      9'b100101011 : begin
        result = input_299;
      end
      9'b100101100 : begin
        result = input_300;
      end
      9'b100101101 : begin
        result = input_301;
      end
      9'b100101110 : begin
        result = input_302;
      end
      9'b100101111 : begin
        result = input_303;
      end
      9'b100110000 : begin
        result = input_304;
      end
      9'b100110001 : begin
        result = input_305;
      end
      9'b100110010 : begin
        result = input_306;
      end
      9'b100110011 : begin
        result = input_307;
      end
      9'b100110100 : begin
        result = input_308;
      end
      9'b100110101 : begin
        result = input_309;
      end
      9'b100110110 : begin
        result = input_310;
      end
      9'b100110111 : begin
        result = input_311;
      end
      9'b100111000 : begin
        result = input_312;
      end
      9'b100111001 : begin
        result = input_313;
      end
      9'b100111010 : begin
        result = input_314;
      end
      9'b100111011 : begin
        result = input_315;
      end
      9'b100111100 : begin
        result = input_316;
      end
      9'b100111101 : begin
        result = input_317;
      end
      9'b100111110 : begin
        result = input_318;
      end
      9'b100111111 : begin
        result = input_319;
      end
      9'b101000000 : begin
        result = input_320;
      end
      9'b101000001 : begin
        result = input_321;
      end
      9'b101000010 : begin
        result = input_322;
      end
      9'b101000011 : begin
        result = input_323;
      end
      9'b101000100 : begin
        result = input_324;
      end
      9'b101000101 : begin
        result = input_325;
      end
      9'b101000110 : begin
        result = input_326;
      end
      9'b101000111 : begin
        result = input_327;
      end
      9'b101001000 : begin
        result = input_328;
      end
      9'b101001001 : begin
        result = input_329;
      end
      9'b101001010 : begin
        result = input_330;
      end
      9'b101001011 : begin
        result = input_331;
      end
      9'b101001100 : begin
        result = input_332;
      end
      9'b101001101 : begin
        result = input_333;
      end
      9'b101001110 : begin
        result = input_334;
      end
      9'b101001111 : begin
        result = input_335;
      end
      9'b101010000 : begin
        result = input_336;
      end
      9'b101010001 : begin
        result = input_337;
      end
      9'b101010010 : begin
        result = input_338;
      end
      9'b101010011 : begin
        result = input_339;
      end
      9'b101010100 : begin
        result = input_340;
      end
      9'b101010101 : begin
        result = input_341;
      end
      9'b101010110 : begin
        result = input_342;
      end
      9'b101010111 : begin
        result = input_343;
      end
      9'b101011000 : begin
        result = input_344;
      end
      9'b101011001 : begin
        result = input_345;
      end
      9'b101011010 : begin
        result = input_346;
      end
      9'b101011011 : begin
        result = input_347;
      end
      9'b101011100 : begin
        result = input_348;
      end
      9'b101011101 : begin
        result = input_349;
      end
      9'b101011110 : begin
        result = input_350;
      end
      9'b101011111 : begin
        result = input_351;
      end
      9'b101100000 : begin
        result = input_352;
      end
      9'b101100001 : begin
        result = input_353;
      end
      9'b101100010 : begin
        result = input_354;
      end
      9'b101100011 : begin
        result = input_355;
      end
      9'b101100100 : begin
        result = input_356;
      end
      9'b101100101 : begin
        result = input_357;
      end
      9'b101100110 : begin
        result = input_358;
      end
      9'b101100111 : begin
        result = input_359;
      end
      9'b101101000 : begin
        result = input_360;
      end
      9'b101101001 : begin
        result = input_361;
      end
      9'b101101010 : begin
        result = input_362;
      end
      9'b101101011 : begin
        result = input_363;
      end
      9'b101101100 : begin
        result = input_364;
      end
      9'b101101101 : begin
        result = input_365;
      end
      9'b101101110 : begin
        result = input_366;
      end
      9'b101101111 : begin
        result = input_367;
      end
      9'b101110000 : begin
        result = input_368;
      end
      9'b101110001 : begin
        result = input_369;
      end
      9'b101110010 : begin
        result = input_370;
      end
      9'b101110011 : begin
        result = input_371;
      end
      9'b101110100 : begin
        result = input_372;
      end
      9'b101110101 : begin
        result = input_373;
      end
      9'b101110110 : begin
        result = input_374;
      end
      9'b101110111 : begin
        result = input_375;
      end
      9'b101111000 : begin
        result = input_376;
      end
      9'b101111001 : begin
        result = input_377;
      end
      9'b101111010 : begin
        result = input_378;
      end
      9'b101111011 : begin
        result = input_379;
      end
      9'b101111100 : begin
        result = input_380;
      end
      9'b101111101 : begin
        result = input_381;
      end
      9'b101111110 : begin
        result = input_382;
      end
      default : begin
        result = input_383;
      end
    endcase
    MUX_v_16_384_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_3_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [1:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_16_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [15:0] readslicef_20_16_4;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_20_16_4 = tmp[15:0];
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_2;
    input [1:0] vector;
  begin
    signext_4_2= {{2{vector[1]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_2_8 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_8 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    myproject
// ------------------------------------------------------------------


module myproject (
  clk, rst, input_1_rsc_dat, layer6_out_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer6_out_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  converterBlock_myproject_core myproject_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .layer6_out_rsc_dat(layer6_out_rsc_dat)
    );
endmodule



