
//------> ./myproject_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module converterBlock_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./myproject_ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module converterBlock_ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./myproject.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
// 
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Thu Oct 27 16:10:15 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core
// ------------------------------------------------------------------


module converterBlock_myproject_core (
  clk, rst, input_1_rsc_dat, layer5_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer5_out_rsc_dat;
  input [8959:0] w2_rsc_dat;
  input [639:0] b2_rsc_dat;
  input [1919:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;


  // Interconnect Declarations
  wire [223:0] input_1_rsci_idat;
  wire [8959:0] w2_rsci_idat;
  wire [639:0] b2_rsci_idat;
  wire [1919:0] w5_rsci_idat;
  wire [14:0] b5_rsci_idat;
  reg [15:0] layer5_out_rsci_idat_47_32;
  wire [21:0] nl_layer5_out_rsci_idat_47_32;
  reg [15:0] layer5_out_rsci_idat_31_16;
  wire [21:0] nl_layer5_out_rsci_idat_31_16;
  reg [15:0] layer5_out_rsci_idat_15_0;
  wire [21:0] nl_layer5_out_rsci_idat_15_0;
  wire [15:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [16:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1;
  wire [15:0] layer2_out_0_sva_1;
  wire [16:0] nl_layer2_out_0_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_0;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_9;
  wire [7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_8_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_0;
  wire layer4_out_conc_193_9;
  wire [7:0] layer4_out_conc_193_8_1;
  wire layer4_out_conc_193_0;
  wire layer4_out_conc_195_9;
  wire [7:0] layer4_out_conc_195_8_1;
  wire layer4_out_conc_195_0;
  wire layer4_out_conc_197_9;
  wire [7:0] layer4_out_conc_197_8_1;
  wire layer4_out_conc_197_0;
  wire layer4_out_conc_199_9;
  wire [7:0] layer4_out_conc_199_8_1;
  wire layer4_out_conc_199_0;
  wire layer4_out_conc_201_9;
  wire [7:0] layer4_out_conc_201_8_1;
  wire layer4_out_conc_201_0;
  wire layer4_out_conc_203_9;
  wire [7:0] layer4_out_conc_203_8_1;
  wire layer4_out_conc_203_0;
  wire layer4_out_conc_205_9;
  wire [7:0] layer4_out_conc_205_8_1;
  wire layer4_out_conc_205_0;
  wire layer4_out_conc_207_9;
  wire [7:0] layer4_out_conc_207_8_1;
  wire layer4_out_conc_207_0;
  wire layer4_out_conc_209_9;
  wire [7:0] layer4_out_conc_209_8_1;
  wire layer4_out_conc_209_0;
  wire layer4_out_conc_211_9;
  wire [7:0] layer4_out_conc_211_8_1;
  wire layer4_out_conc_211_0;
  wire layer4_out_conc_213_9;
  wire [7:0] layer4_out_conc_213_8_1;
  wire layer4_out_conc_213_0;
  wire layer4_out_conc_215_9;
  wire [7:0] layer4_out_conc_215_8_1;
  wire layer4_out_conc_215_0;
  wire layer4_out_conc_217_9;
  wire [7:0] layer4_out_conc_217_8_1;
  wire layer4_out_conc_217_0;
  wire layer4_out_conc_219_9;
  wire [7:0] layer4_out_conc_219_8_1;
  wire layer4_out_conc_219_0;
  wire layer4_out_conc_221_9;
  wire [7:0] layer4_out_conc_221_8_1;
  wire layer4_out_conc_221_0;
  wire layer4_out_conc_223_9;
  wire [7:0] layer4_out_conc_223_8_1;
  wire layer4_out_conc_223_0;
  wire layer4_out_conc_225_9;
  wire [7:0] layer4_out_conc_225_8_1;
  wire layer4_out_conc_225_0;
  wire layer4_out_conc_227_9;
  wire [7:0] layer4_out_conc_227_8_1;
  wire layer4_out_conc_227_0;
  wire layer4_out_conc_229_9;
  wire [7:0] layer4_out_conc_229_8_1;
  wire layer4_out_conc_229_0;
  wire layer4_out_conc_231_9;
  wire [7:0] layer4_out_conc_231_8_1;
  wire layer4_out_conc_231_0;
  wire layer4_out_conc_233_9;
  wire [7:0] layer4_out_conc_233_8_1;
  wire layer4_out_conc_233_0;
  wire layer4_out_conc_235_9;
  wire [7:0] layer4_out_conc_235_8_1;
  wire layer4_out_conc_235_0;
  wire layer4_out_conc_237_9;
  wire [7:0] layer4_out_conc_237_8_1;
  wire layer4_out_conc_237_0;
  wire layer4_out_conc_239_9;
  wire [7:0] layer4_out_conc_239_8_1;
  wire layer4_out_conc_239_0;
  wire layer4_out_conc_241_9;
  wire [7:0] layer4_out_conc_241_8_1;
  wire layer4_out_conc_241_0;
  wire layer4_out_conc_243_9;
  wire [7:0] layer4_out_conc_243_8_1;
  wire layer4_out_conc_243_0;
  wire layer4_out_conc_245_9;
  wire [7:0] layer4_out_conc_245_8_1;
  wire layer4_out_conc_245_0;
  wire layer4_out_conc_247_9;
  wire [7:0] layer4_out_conc_247_8_1;
  wire layer4_out_conc_247_0;
  wire layer4_out_conc_249_9;
  wire [7:0] layer4_out_conc_249_8_1;
  wire layer4_out_conc_249_0;
  wire layer4_out_conc_251_9;
  wire [7:0] layer4_out_conc_251_8_1;
  wire layer4_out_conc_251_0;
  wire layer4_out_conc_253_9;
  wire [7:0] layer4_out_conc_253_8_1;
  wire layer4_out_conc_253_0;
  wire layer4_out_conc_255_9;
  wire [7:0] layer4_out_conc_255_8_1;
  wire layer4_out_conc_255_0;
  wire layer4_out_conc_257_9;
  wire [7:0] layer4_out_conc_257_8_1;
  wire layer4_out_conc_257_0;
  wire layer4_out_conc_259_9;
  wire [7:0] layer4_out_conc_259_8_1;
  wire layer4_out_conc_259_0;
  wire layer4_out_conc_261_9;
  wire [7:0] layer4_out_conc_261_8_1;
  wire layer4_out_conc_261_0;
  wire layer4_out_conc_263_9;
  wire [7:0] layer4_out_conc_263_8_1;
  wire layer4_out_conc_263_0;
  wire layer4_out_conc_265_9;
  wire [7:0] layer4_out_conc_265_8_1;
  wire layer4_out_conc_265_0;
  wire layer4_out_conc_267_9;
  wire [7:0] layer4_out_conc_267_8_1;
  wire layer4_out_conc_267_0;
  wire layer4_out_conc_269_9;
  wire [7:0] layer4_out_conc_269_8_1;
  wire layer4_out_conc_269_0;
  wire layer4_out_conc_271_9;
  wire [7:0] layer4_out_conc_271_8_1;
  wire layer4_out_conc_271_0;
  wire layer4_out_conc_273_9;
  wire [7:0] layer4_out_conc_273_8_1;
  wire layer4_out_conc_273_0;
  wire layer4_out_conc_275_9;
  wire [7:0] layer4_out_conc_275_8_1;
  wire layer4_out_conc_275_0;
  wire layer4_out_conc_277_9;
  wire [7:0] layer4_out_conc_277_8_1;
  wire layer4_out_conc_277_0;
  wire layer4_out_conc_279_9;
  wire [7:0] layer4_out_conc_279_8_1;
  wire layer4_out_conc_279_0;
  wire layer4_out_conc_281_9;
  wire [7:0] layer4_out_conc_281_8_1;
  wire layer4_out_conc_281_0;
  wire layer4_out_conc_283_9;
  wire [7:0] layer4_out_conc_283_8_1;
  wire layer4_out_conc_283_0;
  wire layer4_out_conc_285_9;
  wire [7:0] layer4_out_conc_285_8_1;
  wire layer4_out_conc_285_0;
  wire layer4_out_conc_287_9;
  wire [7:0] layer4_out_conc_287_8_1;
  wire layer4_out_conc_287_0;
  wire layer4_out_conc_289_9;
  wire [7:0] layer4_out_conc_289_8_1;
  wire layer4_out_conc_289_0;
  wire layer4_out_conc_291_9;
  wire [7:0] layer4_out_conc_291_8_1;
  wire layer4_out_conc_291_0;
  wire layer4_out_conc_293_9;
  wire [7:0] layer4_out_conc_293_8_1;
  wire layer4_out_conc_293_0;
  wire layer4_out_conc_295_9;
  wire [7:0] layer4_out_conc_295_8_1;
  wire layer4_out_conc_295_0;
  wire layer4_out_conc_297_9;
  wire [7:0] layer4_out_conc_297_8_1;
  wire layer4_out_conc_297_0;
  wire layer4_out_conc_299_9;
  wire [7:0] layer4_out_conc_299_8_1;
  wire layer4_out_conc_299_0;
  wire layer4_out_conc_301_9;
  wire [7:0] layer4_out_conc_301_8_1;
  wire layer4_out_conc_301_0;
  wire layer4_out_conc_303_9;
  wire [7:0] layer4_out_conc_303_8_1;
  wire layer4_out_conc_303_0;
  wire layer4_out_conc_305_9;
  wire [7:0] layer4_out_conc_305_8_1;
  wire layer4_out_conc_305_0;
  wire layer4_out_conc_307_9;
  wire [7:0] layer4_out_conc_307_8_1;
  wire layer4_out_conc_307_0;
  wire layer4_out_conc_309_9;
  wire [7:0] layer4_out_conc_309_8_1;
  wire layer4_out_conc_309_0;
  wire layer4_out_conc_311_9;
  wire [7:0] layer4_out_conc_311_8_1;
  wire layer4_out_conc_311_0;
  wire layer4_out_conc_313_9;
  wire [7:0] layer4_out_conc_313_8_1;
  wire layer4_out_conc_313_0;
  wire layer4_out_conc_315_9;
  wire [7:0] layer4_out_conc_315_8_1;
  wire layer4_out_conc_315_0;
  wire layer4_out_conc_317_9;
  wire [7:0] layer4_out_conc_317_8_1;
  wire layer4_out_conc_317_0;
  wire layer4_out_conc_319_9;
  wire [7:0] layer4_out_conc_319_8_1;
  wire layer4_out_conc_319_0;
  wire [10:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1;
  wire [10:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1;
  wire [10:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  wire [15:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;
  wire [15:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1;

  wire[15:0] ACCUM_INNER_LOOP_1_acc_393_nl;
  wire[21:0] nl_ACCUM_INNER_LOOP_1_acc_393_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_1_acc_392_nl;
  wire[20:0] nl_ACCUM_INNER_LOOP_1_acc_392_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl;
  wire[5:0] ACCUM_INNER_LOOP_1_acc_396_nl;
  wire[6:0] nl_ACCUM_INNER_LOOP_1_acc_396_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_1_acc_266_nl;
  wire[21:0] nl_ACCUM_INNER_LOOP_1_acc_266_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_1_acc_265_nl;
  wire[20:0] nl_ACCUM_INNER_LOOP_1_acc_265_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl;
  wire[5:0] ACCUM_INNER_LOOP_1_acc_395_nl;
  wire[6:0] nl_ACCUM_INNER_LOOP_1_acc_395_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_1_acc_139_nl;
  wire[21:0] nl_ACCUM_INNER_LOOP_1_acc_139_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_1_acc_140_nl;
  wire[20:0] nl_ACCUM_INNER_LOOP_1_acc_140_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl;
  wire[5:0] ACCUM_INNER_LOOP_1_acc_397_nl;
  wire[6:0] nl_ACCUM_INNER_LOOP_1_acc_397_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_17_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_17_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_13_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_13_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_16_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_16_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1669_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1669_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_30_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_30_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_29_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_29_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_26_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_26_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_25_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_25_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1670_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1670_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_43_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_43_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_42_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_42_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_39_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_39_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_38_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_38_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1671_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1671_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_56_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_56_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_55_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_55_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_52_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_52_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_51_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_51_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1672_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1672_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_69_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_69_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_68_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_68_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_65_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_65_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_64_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_64_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1673_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1673_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_82_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_82_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_81_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_81_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_78_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_78_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_77_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_77_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1674_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1674_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_95_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_95_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_94_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_94_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_91_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_91_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_90_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_90_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1675_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1675_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_108_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_108_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_107_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_107_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_104_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_104_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_103_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_103_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1676_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1676_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_121_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_121_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_120_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_120_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_117_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_117_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_116_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_116_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1677_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1677_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_134_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_134_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_133_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_133_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_130_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_130_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_129_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_129_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1678_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1678_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_147_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_147_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_146_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_146_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_143_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_143_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_142_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_142_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1679_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1679_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_160_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_160_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_159_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_159_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_156_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_156_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_155_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_155_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1680_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1680_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_173_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_173_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_172_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_172_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_169_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_169_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_168_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_168_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1681_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1681_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_186_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_186_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_185_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_185_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_182_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_182_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_181_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_181_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1682_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1682_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_199_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_199_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_198_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_198_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_195_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_195_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_194_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_194_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1683_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1683_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_212_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_212_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_211_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_211_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_208_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_208_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_207_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_207_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1684_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1684_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_225_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_225_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_224_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_224_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_221_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_221_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_220_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_220_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1685_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1685_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_238_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_238_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_237_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_237_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_234_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_234_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_233_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_233_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1686_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1686_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_251_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_251_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_250_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_250_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_247_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_247_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_246_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_246_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1687_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1687_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_264_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_264_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_263_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_263_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_260_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_260_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_259_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_259_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1688_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1688_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_277_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_277_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_276_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_276_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_273_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_273_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_272_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_272_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1689_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1689_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_290_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_290_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_289_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_289_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_286_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_286_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_285_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_285_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1690_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1690_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_303_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_303_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_302_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_302_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_299_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_299_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_298_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_298_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1691_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1691_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_316_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_316_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_315_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_315_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_312_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_312_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_311_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_311_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1692_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1692_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_329_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_329_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_328_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_328_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_325_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_325_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_324_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_324_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1693_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1693_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_342_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_342_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_341_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_341_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_338_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_338_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_337_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_337_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1694_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1694_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_355_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_355_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_354_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_354_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_351_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_351_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_350_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_350_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1695_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1695_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_368_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_368_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_367_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_367_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_364_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_364_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_363_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_363_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1696_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1696_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_381_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_381_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_380_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_380_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_377_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_377_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_376_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_376_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1697_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1697_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_394_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_394_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_393_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_393_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_390_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_390_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_389_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_389_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1698_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1698_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_407_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_407_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_406_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_406_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_403_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_403_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_402_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_402_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1699_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1699_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_420_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_420_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_419_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_419_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_416_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_416_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_415_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_415_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1700_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1700_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_433_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_433_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_432_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_432_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_429_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_429_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_428_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_428_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1701_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1701_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_446_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_446_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_445_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_445_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_442_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_442_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_441_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_441_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1702_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1702_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_459_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_459_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_458_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_458_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_455_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_455_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_454_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_454_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1703_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1703_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_472_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_472_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_471_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_471_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_468_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_468_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_467_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_467_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1704_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1704_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_485_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_485_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_484_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_484_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_481_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_481_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_480_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_480_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1705_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1705_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_498_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_498_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_497_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_497_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_494_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_494_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_493_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_493_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1706_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1706_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_511_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_511_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_510_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_510_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_507_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_507_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_506_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_506_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1707_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1707_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_524_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_524_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_523_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_523_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_520_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_520_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_519_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_519_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1708_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1708_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_537_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_537_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_536_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_536_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_533_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_533_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_532_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_532_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1709_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1709_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_550_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_550_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_549_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_549_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_546_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_546_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_545_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_545_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1710_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1710_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_563_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_563_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_562_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_562_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_559_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_559_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_558_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_558_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1711_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1711_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_576_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_576_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_575_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_575_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_572_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_572_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_571_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_571_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1712_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1712_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_589_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_589_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_588_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_588_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_585_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_585_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_584_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_584_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1713_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1713_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_602_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_602_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_601_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_601_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_598_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_598_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_597_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_597_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1714_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1714_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_615_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_615_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_614_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_614_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_611_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_611_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_610_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_610_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1715_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1715_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_628_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_628_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_627_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_627_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_624_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_624_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_623_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_623_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1716_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1716_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_641_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_641_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_640_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_640_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_637_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_637_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_636_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_636_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1717_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1717_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_654_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_654_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_653_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_653_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_650_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_650_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_649_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_649_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1718_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1718_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_667_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_667_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_666_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_666_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_663_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_663_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_662_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_662_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1719_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1719_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_680_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_680_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_679_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_679_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_676_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_676_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_675_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_675_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1720_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1720_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_693_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_693_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_692_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_692_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_689_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_689_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_688_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_688_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1721_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1721_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_706_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_706_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_705_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_705_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_702_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_702_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_701_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_701_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1722_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1722_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_719_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_719_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_718_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_718_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_715_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_715_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_714_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_714_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1723_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1723_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_732_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_732_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_731_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_731_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_728_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_728_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_727_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_727_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1724_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1724_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_745_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_745_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_744_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_744_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_741_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_741_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_740_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_740_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1725_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1725_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_758_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_758_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_757_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_757_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_754_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_754_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_753_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_753_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1726_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1726_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_771_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_771_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_770_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_770_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_767_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_767_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_766_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_766_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1727_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1727_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_784_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_784_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_783_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_783_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_780_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_780_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_779_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_779_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1728_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1728_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_797_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_797_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_796_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_796_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_793_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_793_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_792_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_792_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1729_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1729_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_810_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_810_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_809_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_809_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_806_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_806_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_805_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_805_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1730_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1730_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_823_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_823_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_822_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_822_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_819_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_819_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_818_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_818_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1731_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1731_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_836_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_836_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_835_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_835_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_832_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_832_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_831_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_831_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1732_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1732_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_849_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_849_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_848_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_848_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_845_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_845_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_844_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_844_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1733_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1733_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_862_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_862_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_861_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_861_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_858_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_858_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_857_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_857_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1734_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1734_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_875_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_875_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_874_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_874_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_871_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_871_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_870_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_870_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1735_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1735_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_888_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_888_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_887_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_887_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_884_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_884_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_883_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_883_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1736_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1736_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_901_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_901_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_900_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_900_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_897_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_897_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_896_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_896_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1737_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1737_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_914_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_914_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_913_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_913_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_910_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_910_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_909_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_909_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1738_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1738_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_927_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_927_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_926_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_926_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_923_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_923_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_922_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_922_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1739_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1739_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_940_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_940_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_939_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_939_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_936_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_936_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_935_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_935_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1740_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1740_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_953_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_953_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_952_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_952_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_949_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_949_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_948_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_948_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1741_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1741_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_966_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_966_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_965_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_965_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_962_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_962_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_961_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_961_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1742_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1742_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_979_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_979_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_978_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_978_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_975_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_975_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_974_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_974_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1743_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1743_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_992_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_992_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_991_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_991_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_988_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_988_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_987_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_987_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1744_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1744_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1005_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1005_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1004_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1004_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1001_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1001_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1000_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1000_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1745_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1745_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1018_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1018_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1017_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1017_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1014_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1014_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1013_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1013_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1746_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1746_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1031_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1031_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1030_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1030_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1027_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1027_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1026_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1026_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1747_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1747_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1044_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1044_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1043_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1043_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1040_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1040_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1039_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1039_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1748_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1748_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1057_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1057_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1056_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1056_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1053_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1053_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1052_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1052_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1749_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1749_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1070_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1070_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1069_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1069_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1066_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1066_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1065_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1065_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1750_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1750_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1083_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1083_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1082_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1082_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1079_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1079_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1078_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1078_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1751_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1751_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1096_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1096_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1095_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1095_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1092_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1092_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1091_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1091_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1752_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1752_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1109_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1109_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1108_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1108_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1105_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1105_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1104_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1104_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1753_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1753_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1122_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1122_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1121_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1121_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1118_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1118_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1117_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1117_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1754_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1754_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1135_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1135_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1134_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1134_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1131_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1131_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1130_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1130_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1755_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1755_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1148_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1148_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1147_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1147_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1144_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1144_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1143_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1143_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1756_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1756_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1161_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1161_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1160_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1160_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1157_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1157_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1156_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1156_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1757_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1757_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1174_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1174_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1173_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1173_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1170_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1170_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1169_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1169_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1758_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1758_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1187_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1187_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1186_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1186_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1183_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1183_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1182_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1182_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1759_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1759_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1200_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1200_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1199_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1199_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1196_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1196_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1195_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1195_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1760_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1760_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1213_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1213_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1212_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1212_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1209_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1209_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1208_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1208_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1761_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1761_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1226_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1226_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1225_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1225_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1222_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1222_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1221_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1221_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1762_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1762_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1239_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1239_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1238_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1238_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1235_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1235_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1234_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1234_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1763_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1763_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1252_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1252_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1251_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1251_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1248_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1248_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1247_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1247_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1764_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1764_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1265_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1265_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1264_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1264_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1261_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1261_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1260_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1260_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1765_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1765_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1278_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1278_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1277_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1277_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1274_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1274_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1273_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1273_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1766_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1766_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1291_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1291_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1290_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1290_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1287_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1287_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1286_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1286_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1767_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1767_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1304_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1304_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1303_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1303_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1300_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1300_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1299_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1299_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1768_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1768_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1317_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1317_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1316_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1316_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1313_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1313_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1312_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1312_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1769_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1769_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1330_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1330_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1329_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1329_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1326_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1326_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1325_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1325_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1770_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1770_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1343_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1343_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1342_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1342_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1339_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1339_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1338_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1338_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1771_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1771_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1356_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1356_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1355_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1355_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1352_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1352_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1351_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1351_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1772_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1772_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1369_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1369_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1368_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1368_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1365_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1365_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1364_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1364_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1773_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1773_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1382_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1382_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1381_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1381_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1378_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1378_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1377_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1377_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1774_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1774_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1395_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1395_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1394_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1394_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1391_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1391_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1390_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1390_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1775_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1775_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1408_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1408_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1407_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1407_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1404_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1404_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1403_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1403_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1776_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1776_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1421_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1421_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1420_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1420_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1417_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1417_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1416_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1416_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1777_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1777_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1434_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1434_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1433_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1433_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1430_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1430_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1429_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1429_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1778_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1778_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1447_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1447_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1446_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1446_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1443_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1443_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1442_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1442_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1779_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1779_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1460_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1460_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1459_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1459_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1456_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1456_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1455_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1455_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1780_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1780_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1473_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1473_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1472_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1472_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1469_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1469_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1468_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1468_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1781_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1781_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1486_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1486_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1485_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1485_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1482_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1482_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1481_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1481_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1782_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1782_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1499_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1499_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1498_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1498_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1495_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1495_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1494_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1494_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1783_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1783_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1512_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1512_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1511_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1511_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1508_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1508_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1507_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1507_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1784_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1784_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1525_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1525_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1524_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1524_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1521_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1521_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1520_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1520_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1785_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1785_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1538_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1538_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1537_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1537_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1534_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1534_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1533_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1533_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1786_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1786_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1551_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1551_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1550_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1550_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1547_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1547_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1546_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1546_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1787_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1787_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1564_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1564_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1563_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1563_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1560_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1560_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1559_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1559_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1788_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1788_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1577_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1577_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1576_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1576_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1573_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1573_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1572_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1572_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1789_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1789_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1590_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1590_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1589_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1589_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1586_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1586_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1585_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1585_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1790_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1790_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1603_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1603_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1602_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1602_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1599_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1599_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1598_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1598_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1791_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1791_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1616_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1616_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1615_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1615_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1612_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1612_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1611_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1611_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1792_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1792_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1629_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1629_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1628_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1628_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1625_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1625_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1624_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1624_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1793_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1793_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1642_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1642_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1641_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1641_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1638_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1638_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1637_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1637_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1794_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1794_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1655_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1655_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1654_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1654_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1651_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1651_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1650_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1650_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1795_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1795_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1668_nl;
  wire[18:0] nl_ACCUM_INNER_LOOP_acc_1668_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1667_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1667_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1664_nl;
  wire[17:0] nl_ACCUM_INNER_LOOP_acc_1664_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl;
  wire[15:0] ACCUM_INNER_LOOP_acc_1663_nl;
  wire[16:0] nl_ACCUM_INNER_LOOP_acc_1663_nl;
  wire[9:0] ACCUM_INNER_LOOP_acc_1796_nl;
  wire[10:0] nl_ACCUM_INNER_LOOP_acc_1796_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl;
  wire[14:0] ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl;
  wire signed [15:0] nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[16:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[19:0] ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire signed [20:0] nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;
  wire[7:0] nnet_relu_layer2_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [47:0] nl_layer5_out_rsci_idat;
  assign nl_layer5_out_rsci_idat = {layer5_out_rsci_idat_47_32 , layer5_out_rsci_idat_31_16
      , layer5_out_rsci_idat_15_0};
  converterBlock_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd224)) input_1_rsci (
      .dat(input_1_rsc_dat),
      .idat(input_1_rsci_idat)
    );
  converterBlock_ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd48)) layer5_out_rsci (
      .idat(nl_layer5_out_rsci_idat[47:0]),
      .dat(layer5_out_rsc_dat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd8960)) w2_rsci (
      .dat(w2_rsc_dat),
      .idat(w2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd640)) b2_rsci (
      .dat(b2_rsc_dat),
      .idat(b2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd1920)) w5_rsci (
      .dat(w5_rsc_dat),
      .idat(w5_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd15)) b5_rsci (
      .dat(b5_rsc_dat),
      .idat(b5_rsci_idat)
    );
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1 = (layer2_out_0_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[29:25]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[34:30]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[9:5]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[14:10]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[19:15]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[24:20]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[39:35]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[44:40]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_17_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_17_nl = nl_ACCUM_INNER_LOOP_acc_17_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[49:45]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[54:50]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[59:55]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[64:60]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_13_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_13_nl = nl_ACCUM_INNER_LOOP_acc_13_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1669_nl = (ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[4:0]);
  assign ACCUM_INNER_LOOP_acc_1669_nl = nl_ACCUM_INNER_LOOP_acc_1669_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4:0]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_16_nl = ({ACCUM_INNER_LOOP_acc_1669_nl , (ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_16_nl = nl_ACCUM_INNER_LOOP_acc_16_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_nl = ACCUM_INNER_LOOP_acc_13_nl + ACCUM_INNER_LOOP_acc_16_nl;
  assign ACCUM_INNER_LOOP_acc_nl = nl_ACCUM_INNER_LOOP_acc_nl[15:0];
  assign nl_layer2_out_0_sva_1 = ACCUM_INNER_LOOP_acc_17_nl + ACCUM_INNER_LOOP_acc_nl;
  assign layer2_out_0_sva_1 = nl_layer2_out_0_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 = (ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[99:95]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[104:100]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[79:75]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[84:80]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[89:85]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[94:90]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[109:105]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[114:110]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_30_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_30_nl = nl_ACCUM_INNER_LOOP_acc_30_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[119:115]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[124:120]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[129:125]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[134:130]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_26_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_26_nl = nl_ACCUM_INNER_LOOP_acc_26_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1670_nl = (ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[9:5]);
  assign ACCUM_INNER_LOOP_acc_1670_nl = nl_ACCUM_INNER_LOOP_acc_1670_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[74:70]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_25_nl = ({ACCUM_INNER_LOOP_acc_1670_nl , (ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_25_nl = nl_ACCUM_INNER_LOOP_acc_25_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_29_nl = ACCUM_INNER_LOOP_acc_26_nl + ACCUM_INNER_LOOP_acc_25_nl;
  assign ACCUM_INNER_LOOP_acc_29_nl = nl_ACCUM_INNER_LOOP_acc_29_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_30_nl
      + ACCUM_INNER_LOOP_acc_29_nl;
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 = (ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[169:165]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[174:170]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[149:145]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[154:150]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[159:155]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[164:160]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[179:175]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[184:180]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_43_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_43_nl = nl_ACCUM_INNER_LOOP_acc_43_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[189:185]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[194:190]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[199:195]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[204:200]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_39_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_39_nl = nl_ACCUM_INNER_LOOP_acc_39_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1671_nl = (ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[14:10]);
  assign ACCUM_INNER_LOOP_acc_1671_nl = nl_ACCUM_INNER_LOOP_acc_1671_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[144:140]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_38_nl = ({ACCUM_INNER_LOOP_acc_1671_nl , (ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_38_nl = nl_ACCUM_INNER_LOOP_acc_38_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_42_nl = ACCUM_INNER_LOOP_acc_39_nl + ACCUM_INNER_LOOP_acc_38_nl;
  assign ACCUM_INNER_LOOP_acc_42_nl = nl_ACCUM_INNER_LOOP_acc_42_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_43_nl
      + ACCUM_INNER_LOOP_acc_42_nl;
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 = (ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[239:235]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[244:240]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[219:215]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[224:220]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[229:225]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[234:230]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[249:245]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[254:250]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_56_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_56_nl = nl_ACCUM_INNER_LOOP_acc_56_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[259:255]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[264:260]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[269:265]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[274:270]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_52_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_52_nl = nl_ACCUM_INNER_LOOP_acc_52_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1672_nl = (ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[19:15]);
  assign ACCUM_INNER_LOOP_acc_1672_nl = nl_ACCUM_INNER_LOOP_acc_1672_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[214:210]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_51_nl = ({ACCUM_INNER_LOOP_acc_1672_nl , (ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_51_nl = nl_ACCUM_INNER_LOOP_acc_51_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_55_nl = ACCUM_INNER_LOOP_acc_52_nl + ACCUM_INNER_LOOP_acc_51_nl;
  assign ACCUM_INNER_LOOP_acc_55_nl = nl_ACCUM_INNER_LOOP_acc_55_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_56_nl
      + ACCUM_INNER_LOOP_acc_55_nl;
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 = (ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[309:305]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[314:310]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[289:285]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[294:290]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[299:295]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[304:300]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[319:315]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[324:320]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_69_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_69_nl = nl_ACCUM_INNER_LOOP_acc_69_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[329:325]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[334:330]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[339:335]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[344:340]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_65_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_65_nl = nl_ACCUM_INNER_LOOP_acc_65_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1673_nl = (ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[24:20]);
  assign ACCUM_INNER_LOOP_acc_1673_nl = nl_ACCUM_INNER_LOOP_acc_1673_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[284:280]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_64_nl = ({ACCUM_INNER_LOOP_acc_1673_nl , (ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_64_nl = nl_ACCUM_INNER_LOOP_acc_64_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_68_nl = ACCUM_INNER_LOOP_acc_65_nl + ACCUM_INNER_LOOP_acc_64_nl;
  assign ACCUM_INNER_LOOP_acc_68_nl = nl_ACCUM_INNER_LOOP_acc_68_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_69_nl
      + ACCUM_INNER_LOOP_acc_68_nl;
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 = (ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[379:375]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[384:380]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[359:355]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[364:360]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[369:365]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[374:370]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[389:385]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[394:390]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_82_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_82_nl = nl_ACCUM_INNER_LOOP_acc_82_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[399:395]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[404:400]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[409:405]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[414:410]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_78_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_78_nl = nl_ACCUM_INNER_LOOP_acc_78_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1674_nl = (ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[29:25]);
  assign ACCUM_INNER_LOOP_acc_1674_nl = nl_ACCUM_INNER_LOOP_acc_1674_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[354:350]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_77_nl = ({ACCUM_INNER_LOOP_acc_1674_nl , (ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_77_nl = nl_ACCUM_INNER_LOOP_acc_77_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_81_nl = ACCUM_INNER_LOOP_acc_78_nl + ACCUM_INNER_LOOP_acc_77_nl;
  assign ACCUM_INNER_LOOP_acc_81_nl = nl_ACCUM_INNER_LOOP_acc_81_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_82_nl
      + ACCUM_INNER_LOOP_acc_81_nl;
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 = (ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[449:445]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[454:450]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[429:425]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[434:430]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[439:435]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[444:440]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[459:455]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[464:460]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_95_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_95_nl = nl_ACCUM_INNER_LOOP_acc_95_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[469:465]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[474:470]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[479:475]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[484:480]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_91_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_91_nl = nl_ACCUM_INNER_LOOP_acc_91_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1675_nl = (ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[34:30]);
  assign ACCUM_INNER_LOOP_acc_1675_nl = nl_ACCUM_INNER_LOOP_acc_1675_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[424:420]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_90_nl = ({ACCUM_INNER_LOOP_acc_1675_nl , (ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_90_nl = nl_ACCUM_INNER_LOOP_acc_90_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_94_nl = ACCUM_INNER_LOOP_acc_91_nl + ACCUM_INNER_LOOP_acc_90_nl;
  assign ACCUM_INNER_LOOP_acc_94_nl = nl_ACCUM_INNER_LOOP_acc_94_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_95_nl
      + ACCUM_INNER_LOOP_acc_94_nl;
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 = (ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[519:515]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[524:520]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[499:495]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[504:500]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[509:505]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[514:510]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[529:525]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[534:530]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_108_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_108_nl = nl_ACCUM_INNER_LOOP_acc_108_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[539:535]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[544:540]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[549:545]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[554:550]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_104_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_104_nl = nl_ACCUM_INNER_LOOP_acc_104_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1676_nl = (ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[39:35]);
  assign ACCUM_INNER_LOOP_acc_1676_nl = nl_ACCUM_INNER_LOOP_acc_1676_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[494:490]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_103_nl = ({ACCUM_INNER_LOOP_acc_1676_nl , (ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_103_nl = nl_ACCUM_INNER_LOOP_acc_103_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_107_nl = ACCUM_INNER_LOOP_acc_104_nl + ACCUM_INNER_LOOP_acc_103_nl;
  assign ACCUM_INNER_LOOP_acc_107_nl = nl_ACCUM_INNER_LOOP_acc_107_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_108_nl
      + ACCUM_INNER_LOOP_acc_107_nl;
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 = (ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[589:585]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[594:590]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[569:565]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[574:570]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[579:575]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[584:580]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[599:595]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[604:600]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_121_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_121_nl = nl_ACCUM_INNER_LOOP_acc_121_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[609:605]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[614:610]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[619:615]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[624:620]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_117_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_117_nl = nl_ACCUM_INNER_LOOP_acc_117_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1677_nl = (ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[44:40]);
  assign ACCUM_INNER_LOOP_acc_1677_nl = nl_ACCUM_INNER_LOOP_acc_1677_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[564:560]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_116_nl = ({ACCUM_INNER_LOOP_acc_1677_nl , (ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_116_nl = nl_ACCUM_INNER_LOOP_acc_116_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_120_nl = ACCUM_INNER_LOOP_acc_117_nl + ACCUM_INNER_LOOP_acc_116_nl;
  assign ACCUM_INNER_LOOP_acc_120_nl = nl_ACCUM_INNER_LOOP_acc_120_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_121_nl
      + ACCUM_INNER_LOOP_acc_120_nl;
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 = (ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[659:655]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[664:660]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[639:635]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[644:640]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[649:645]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[654:650]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[669:665]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[674:670]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_134_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_134_nl = nl_ACCUM_INNER_LOOP_acc_134_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[679:675]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[684:680]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[689:685]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[694:690]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_130_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_130_nl = nl_ACCUM_INNER_LOOP_acc_130_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1678_nl = (ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[49:45]);
  assign ACCUM_INNER_LOOP_acc_1678_nl = nl_ACCUM_INNER_LOOP_acc_1678_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[634:630]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_129_nl = ({ACCUM_INNER_LOOP_acc_1678_nl , (ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_129_nl = nl_ACCUM_INNER_LOOP_acc_129_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_133_nl = ACCUM_INNER_LOOP_acc_130_nl + ACCUM_INNER_LOOP_acc_129_nl;
  assign ACCUM_INNER_LOOP_acc_133_nl = nl_ACCUM_INNER_LOOP_acc_133_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_134_nl
      + ACCUM_INNER_LOOP_acc_133_nl;
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 = (ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[729:725]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[734:730]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[709:705]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[714:710]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[719:715]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[724:720]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[739:735]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[744:740]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_147_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_147_nl = nl_ACCUM_INNER_LOOP_acc_147_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[749:745]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[754:750]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[759:755]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[764:760]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_143_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_143_nl = nl_ACCUM_INNER_LOOP_acc_143_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1679_nl = (ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[54:50]);
  assign ACCUM_INNER_LOOP_acc_1679_nl = nl_ACCUM_INNER_LOOP_acc_1679_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[704:700]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_142_nl = ({ACCUM_INNER_LOOP_acc_1679_nl , (ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_142_nl = nl_ACCUM_INNER_LOOP_acc_142_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_146_nl = ACCUM_INNER_LOOP_acc_143_nl + ACCUM_INNER_LOOP_acc_142_nl;
  assign ACCUM_INNER_LOOP_acc_146_nl = nl_ACCUM_INNER_LOOP_acc_146_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_147_nl
      + ACCUM_INNER_LOOP_acc_146_nl;
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 = (ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[799:795]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[804:800]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[779:775]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[784:780]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[789:785]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[794:790]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[809:805]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[814:810]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_160_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_160_nl = nl_ACCUM_INNER_LOOP_acc_160_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[819:815]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[824:820]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[829:825]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[834:830]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_156_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_156_nl = nl_ACCUM_INNER_LOOP_acc_156_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1680_nl = (ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[59:55]);
  assign ACCUM_INNER_LOOP_acc_1680_nl = nl_ACCUM_INNER_LOOP_acc_1680_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[774:770]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_155_nl = ({ACCUM_INNER_LOOP_acc_1680_nl , (ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_155_nl = nl_ACCUM_INNER_LOOP_acc_155_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_159_nl = ACCUM_INNER_LOOP_acc_156_nl + ACCUM_INNER_LOOP_acc_155_nl;
  assign ACCUM_INNER_LOOP_acc_159_nl = nl_ACCUM_INNER_LOOP_acc_159_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_160_nl
      + ACCUM_INNER_LOOP_acc_159_nl;
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 = (ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[869:865]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[874:870]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[849:845]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[854:850]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[859:855]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[864:860]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[879:875]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[884:880]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_173_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_173_nl = nl_ACCUM_INNER_LOOP_acc_173_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[889:885]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[894:890]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[899:895]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[904:900]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_169_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_169_nl = nl_ACCUM_INNER_LOOP_acc_169_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1681_nl = (ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[64:60]);
  assign ACCUM_INNER_LOOP_acc_1681_nl = nl_ACCUM_INNER_LOOP_acc_1681_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[844:840]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_168_nl = ({ACCUM_INNER_LOOP_acc_1681_nl , (ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_168_nl = nl_ACCUM_INNER_LOOP_acc_168_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_172_nl = ACCUM_INNER_LOOP_acc_169_nl + ACCUM_INNER_LOOP_acc_168_nl;
  assign ACCUM_INNER_LOOP_acc_172_nl = nl_ACCUM_INNER_LOOP_acc_172_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_173_nl
      + ACCUM_INNER_LOOP_acc_172_nl;
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 = (ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[939:935]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[944:940]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[919:915]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[924:920]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[929:925]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[934:930]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[949:945]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[954:950]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_186_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_186_nl = nl_ACCUM_INNER_LOOP_acc_186_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[959:955]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[964:960]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[969:965]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[974:970]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_182_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_182_nl = nl_ACCUM_INNER_LOOP_acc_182_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1682_nl = (ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[69:65]);
  assign ACCUM_INNER_LOOP_acc_1682_nl = nl_ACCUM_INNER_LOOP_acc_1682_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[914:910]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_181_nl = ({ACCUM_INNER_LOOP_acc_1682_nl , (ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_181_nl = nl_ACCUM_INNER_LOOP_acc_181_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_185_nl = ACCUM_INNER_LOOP_acc_182_nl + ACCUM_INNER_LOOP_acc_181_nl;
  assign ACCUM_INNER_LOOP_acc_185_nl = nl_ACCUM_INNER_LOOP_acc_185_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_186_nl
      + ACCUM_INNER_LOOP_acc_185_nl;
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 = (ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1009:1005]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1014:1010]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[989:985]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[994:990]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[999:995]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1004:1000]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1019:1015]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1024:1020]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_199_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_199_nl = nl_ACCUM_INNER_LOOP_acc_199_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1029:1025]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1034:1030]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1039:1035]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1044:1040]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_195_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_195_nl = nl_ACCUM_INNER_LOOP_acc_195_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1683_nl = (ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[74:70]);
  assign ACCUM_INNER_LOOP_acc_1683_nl = nl_ACCUM_INNER_LOOP_acc_1683_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[984:980]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_194_nl = ({ACCUM_INNER_LOOP_acc_1683_nl , (ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_194_nl = nl_ACCUM_INNER_LOOP_acc_194_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_198_nl = ACCUM_INNER_LOOP_acc_195_nl + ACCUM_INNER_LOOP_acc_194_nl;
  assign ACCUM_INNER_LOOP_acc_198_nl = nl_ACCUM_INNER_LOOP_acc_198_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_199_nl
      + ACCUM_INNER_LOOP_acc_198_nl;
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 = (ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1079:1075]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1084:1080]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1059:1055]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1064:1060]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1069:1065]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1074:1070]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1089:1085]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1094:1090]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_212_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_212_nl = nl_ACCUM_INNER_LOOP_acc_212_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1099:1095]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1104:1100]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1109:1105]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1114:1110]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_208_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_208_nl = nl_ACCUM_INNER_LOOP_acc_208_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1684_nl = (ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[79:75]);
  assign ACCUM_INNER_LOOP_acc_1684_nl = nl_ACCUM_INNER_LOOP_acc_1684_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1054:1050]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_207_nl = ({ACCUM_INNER_LOOP_acc_1684_nl , (ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_207_nl = nl_ACCUM_INNER_LOOP_acc_207_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_211_nl = ACCUM_INNER_LOOP_acc_208_nl + ACCUM_INNER_LOOP_acc_207_nl;
  assign ACCUM_INNER_LOOP_acc_211_nl = nl_ACCUM_INNER_LOOP_acc_211_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_212_nl
      + ACCUM_INNER_LOOP_acc_211_nl;
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 = (ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1149:1145]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1154:1150]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1129:1125]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1134:1130]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1139:1135]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1144:1140]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1159:1155]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1164:1160]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_225_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_225_nl = nl_ACCUM_INNER_LOOP_acc_225_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1169:1165]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1174:1170]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1179:1175]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1184:1180]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_221_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_221_nl = nl_ACCUM_INNER_LOOP_acc_221_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1685_nl = (ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[84:80]);
  assign ACCUM_INNER_LOOP_acc_1685_nl = nl_ACCUM_INNER_LOOP_acc_1685_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1124:1120]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_220_nl = ({ACCUM_INNER_LOOP_acc_1685_nl , (ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_220_nl = nl_ACCUM_INNER_LOOP_acc_220_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_224_nl = ACCUM_INNER_LOOP_acc_221_nl + ACCUM_INNER_LOOP_acc_220_nl;
  assign ACCUM_INNER_LOOP_acc_224_nl = nl_ACCUM_INNER_LOOP_acc_224_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_225_nl
      + ACCUM_INNER_LOOP_acc_224_nl;
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 = (ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1219:1215]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1224:1220]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1199:1195]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1204:1200]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1209:1205]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1214:1210]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1229:1225]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1234:1230]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_238_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_238_nl = nl_ACCUM_INNER_LOOP_acc_238_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1239:1235]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1244:1240]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1249:1245]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1254:1250]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_234_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_234_nl = nl_ACCUM_INNER_LOOP_acc_234_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1686_nl = (ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[89:85]);
  assign ACCUM_INNER_LOOP_acc_1686_nl = nl_ACCUM_INNER_LOOP_acc_1686_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1194:1190]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_233_nl = ({ACCUM_INNER_LOOP_acc_1686_nl , (ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_233_nl = nl_ACCUM_INNER_LOOP_acc_233_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_237_nl = ACCUM_INNER_LOOP_acc_234_nl + ACCUM_INNER_LOOP_acc_233_nl;
  assign ACCUM_INNER_LOOP_acc_237_nl = nl_ACCUM_INNER_LOOP_acc_237_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_238_nl
      + ACCUM_INNER_LOOP_acc_237_nl;
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 = (ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1289:1285]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1294:1290]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1269:1265]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1274:1270]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1279:1275]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1284:1280]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1299:1295]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1304:1300]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_251_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_251_nl = nl_ACCUM_INNER_LOOP_acc_251_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1309:1305]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1314:1310]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1319:1315]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1324:1320]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_247_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_247_nl = nl_ACCUM_INNER_LOOP_acc_247_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1687_nl = (ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[94:90]);
  assign ACCUM_INNER_LOOP_acc_1687_nl = nl_ACCUM_INNER_LOOP_acc_1687_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1264:1260]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_246_nl = ({ACCUM_INNER_LOOP_acc_1687_nl , (ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_246_nl = nl_ACCUM_INNER_LOOP_acc_246_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_250_nl = ACCUM_INNER_LOOP_acc_247_nl + ACCUM_INNER_LOOP_acc_246_nl;
  assign ACCUM_INNER_LOOP_acc_250_nl = nl_ACCUM_INNER_LOOP_acc_250_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_251_nl
      + ACCUM_INNER_LOOP_acc_250_nl;
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 = (ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1359:1355]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1364:1360]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1339:1335]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1344:1340]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1349:1345]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1354:1350]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1369:1365]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1374:1370]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_264_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_264_nl = nl_ACCUM_INNER_LOOP_acc_264_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1379:1375]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1384:1380]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1389:1385]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1394:1390]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_260_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_260_nl = nl_ACCUM_INNER_LOOP_acc_260_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1688_nl = (ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[99:95]);
  assign ACCUM_INNER_LOOP_acc_1688_nl = nl_ACCUM_INNER_LOOP_acc_1688_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1334:1330]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_259_nl = ({ACCUM_INNER_LOOP_acc_1688_nl , (ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_259_nl = nl_ACCUM_INNER_LOOP_acc_259_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_263_nl = ACCUM_INNER_LOOP_acc_260_nl + ACCUM_INNER_LOOP_acc_259_nl;
  assign ACCUM_INNER_LOOP_acc_263_nl = nl_ACCUM_INNER_LOOP_acc_263_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_264_nl
      + ACCUM_INNER_LOOP_acc_263_nl;
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 = (ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1429:1425]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1434:1430]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1409:1405]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1414:1410]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1419:1415]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1424:1420]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1439:1435]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1444:1440]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_277_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_277_nl = nl_ACCUM_INNER_LOOP_acc_277_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1449:1445]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1454:1450]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1459:1455]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1464:1460]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_273_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_273_nl = nl_ACCUM_INNER_LOOP_acc_273_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1689_nl = (ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[104:100]);
  assign ACCUM_INNER_LOOP_acc_1689_nl = nl_ACCUM_INNER_LOOP_acc_1689_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1404:1400]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_272_nl = ({ACCUM_INNER_LOOP_acc_1689_nl , (ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_272_nl = nl_ACCUM_INNER_LOOP_acc_272_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_276_nl = ACCUM_INNER_LOOP_acc_273_nl + ACCUM_INNER_LOOP_acc_272_nl;
  assign ACCUM_INNER_LOOP_acc_276_nl = nl_ACCUM_INNER_LOOP_acc_276_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_277_nl
      + ACCUM_INNER_LOOP_acc_276_nl;
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 = (ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1499:1495]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1504:1500]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1479:1475]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1484:1480]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1489:1485]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1494:1490]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1509:1505]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1514:1510]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_290_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_290_nl = nl_ACCUM_INNER_LOOP_acc_290_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1519:1515]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1524:1520]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1529:1525]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1534:1530]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_286_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_286_nl = nl_ACCUM_INNER_LOOP_acc_286_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1690_nl = (ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[109:105]);
  assign ACCUM_INNER_LOOP_acc_1690_nl = nl_ACCUM_INNER_LOOP_acc_1690_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1474:1470]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_285_nl = ({ACCUM_INNER_LOOP_acc_1690_nl , (ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_285_nl = nl_ACCUM_INNER_LOOP_acc_285_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_289_nl = ACCUM_INNER_LOOP_acc_286_nl + ACCUM_INNER_LOOP_acc_285_nl;
  assign ACCUM_INNER_LOOP_acc_289_nl = nl_ACCUM_INNER_LOOP_acc_289_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_290_nl
      + ACCUM_INNER_LOOP_acc_289_nl;
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 = (ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1569:1565]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1574:1570]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1549:1545]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1554:1550]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1559:1555]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1564:1560]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1579:1575]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1584:1580]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_303_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_303_nl = nl_ACCUM_INNER_LOOP_acc_303_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1589:1585]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1594:1590]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1599:1595]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1604:1600]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_299_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_299_nl = nl_ACCUM_INNER_LOOP_acc_299_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1691_nl = (ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[114:110]);
  assign ACCUM_INNER_LOOP_acc_1691_nl = nl_ACCUM_INNER_LOOP_acc_1691_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1544:1540]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_298_nl = ({ACCUM_INNER_LOOP_acc_1691_nl , (ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_298_nl = nl_ACCUM_INNER_LOOP_acc_298_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_302_nl = ACCUM_INNER_LOOP_acc_299_nl + ACCUM_INNER_LOOP_acc_298_nl;
  assign ACCUM_INNER_LOOP_acc_302_nl = nl_ACCUM_INNER_LOOP_acc_302_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_303_nl
      + ACCUM_INNER_LOOP_acc_302_nl;
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 = (ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1639:1635]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1644:1640]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1619:1615]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1624:1620]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1629:1625]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1634:1630]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1649:1645]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1654:1650]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_316_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_316_nl = nl_ACCUM_INNER_LOOP_acc_316_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1659:1655]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1664:1660]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1669:1665]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1674:1670]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_312_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_312_nl = nl_ACCUM_INNER_LOOP_acc_312_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1692_nl = (ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[119:115]);
  assign ACCUM_INNER_LOOP_acc_1692_nl = nl_ACCUM_INNER_LOOP_acc_1692_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1614:1610]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_311_nl = ({ACCUM_INNER_LOOP_acc_1692_nl , (ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_311_nl = nl_ACCUM_INNER_LOOP_acc_311_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_315_nl = ACCUM_INNER_LOOP_acc_312_nl + ACCUM_INNER_LOOP_acc_311_nl;
  assign ACCUM_INNER_LOOP_acc_315_nl = nl_ACCUM_INNER_LOOP_acc_315_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_316_nl
      + ACCUM_INNER_LOOP_acc_315_nl;
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 = (ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1709:1705]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1714:1710]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1689:1685]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1694:1690]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1699:1695]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1704:1700]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1719:1715]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1724:1720]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_329_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_329_nl = nl_ACCUM_INNER_LOOP_acc_329_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1729:1725]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1734:1730]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1739:1735]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1744:1740]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_325_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_325_nl = nl_ACCUM_INNER_LOOP_acc_325_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1693_nl = (ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[124:120]);
  assign ACCUM_INNER_LOOP_acc_1693_nl = nl_ACCUM_INNER_LOOP_acc_1693_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1684:1680]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_324_nl = ({ACCUM_INNER_LOOP_acc_1693_nl , (ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_324_nl = nl_ACCUM_INNER_LOOP_acc_324_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_328_nl = ACCUM_INNER_LOOP_acc_325_nl + ACCUM_INNER_LOOP_acc_324_nl;
  assign ACCUM_INNER_LOOP_acc_328_nl = nl_ACCUM_INNER_LOOP_acc_328_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_329_nl
      + ACCUM_INNER_LOOP_acc_328_nl;
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 = (ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1779:1775]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1784:1780]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1759:1755]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1764:1760]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1769:1765]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1774:1770]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1789:1785]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1794:1790]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_342_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_342_nl = nl_ACCUM_INNER_LOOP_acc_342_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1799:1795]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1804:1800]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1809:1805]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1814:1810]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_338_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_338_nl = nl_ACCUM_INNER_LOOP_acc_338_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1694_nl = (ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[129:125]);
  assign ACCUM_INNER_LOOP_acc_1694_nl = nl_ACCUM_INNER_LOOP_acc_1694_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1754:1750]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_337_nl = ({ACCUM_INNER_LOOP_acc_1694_nl , (ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_337_nl = nl_ACCUM_INNER_LOOP_acc_337_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_341_nl = ACCUM_INNER_LOOP_acc_338_nl + ACCUM_INNER_LOOP_acc_337_nl;
  assign ACCUM_INNER_LOOP_acc_341_nl = nl_ACCUM_INNER_LOOP_acc_341_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_342_nl
      + ACCUM_INNER_LOOP_acc_341_nl;
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 = (ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1849:1845]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1854:1850]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1829:1825]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1834:1830]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1839:1835]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1844:1840]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1859:1855]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1864:1860]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_355_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_355_nl = nl_ACCUM_INNER_LOOP_acc_355_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1869:1865]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1874:1870]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1879:1875]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1884:1880]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_351_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_351_nl = nl_ACCUM_INNER_LOOP_acc_351_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1695_nl = (ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[134:130]);
  assign ACCUM_INNER_LOOP_acc_1695_nl = nl_ACCUM_INNER_LOOP_acc_1695_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1824:1820]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_350_nl = ({ACCUM_INNER_LOOP_acc_1695_nl , (ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_350_nl = nl_ACCUM_INNER_LOOP_acc_350_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_354_nl = ACCUM_INNER_LOOP_acc_351_nl + ACCUM_INNER_LOOP_acc_350_nl;
  assign ACCUM_INNER_LOOP_acc_354_nl = nl_ACCUM_INNER_LOOP_acc_354_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_355_nl
      + ACCUM_INNER_LOOP_acc_354_nl;
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 = (ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1919:1915]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1924:1920]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1899:1895]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1904:1900]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1909:1905]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1914:1910]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1929:1925]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[1934:1930]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_368_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_368_nl = nl_ACCUM_INNER_LOOP_acc_368_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[1939:1935]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[1944:1940]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[1949:1945]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[1954:1950]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_364_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_364_nl = nl_ACCUM_INNER_LOOP_acc_364_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1696_nl = (ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[139:135]);
  assign ACCUM_INNER_LOOP_acc_1696_nl = nl_ACCUM_INNER_LOOP_acc_1696_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1894:1890]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_363_nl = ({ACCUM_INNER_LOOP_acc_1696_nl , (ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_363_nl = nl_ACCUM_INNER_LOOP_acc_363_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_367_nl = ACCUM_INNER_LOOP_acc_364_nl + ACCUM_INNER_LOOP_acc_363_nl;
  assign ACCUM_INNER_LOOP_acc_367_nl = nl_ACCUM_INNER_LOOP_acc_367_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_368_nl
      + ACCUM_INNER_LOOP_acc_367_nl;
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 = (ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[1989:1985]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[1994:1990]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[1969:1965]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[1974:1970]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[1979:1975]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[1984:1980]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[1999:1995]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2004:2000]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_381_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_381_nl = nl_ACCUM_INNER_LOOP_acc_381_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2009:2005]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2014:2010]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2019:2015]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2024:2020]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_377_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_377_nl = nl_ACCUM_INNER_LOOP_acc_377_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1697_nl = (ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[144:140]);
  assign ACCUM_INNER_LOOP_acc_1697_nl = nl_ACCUM_INNER_LOOP_acc_1697_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[1964:1960]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_376_nl = ({ACCUM_INNER_LOOP_acc_1697_nl , (ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_376_nl = nl_ACCUM_INNER_LOOP_acc_376_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_380_nl = ACCUM_INNER_LOOP_acc_377_nl + ACCUM_INNER_LOOP_acc_376_nl;
  assign ACCUM_INNER_LOOP_acc_380_nl = nl_ACCUM_INNER_LOOP_acc_380_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_381_nl
      + ACCUM_INNER_LOOP_acc_380_nl;
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 = (ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2059:2055]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2064:2060]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2039:2035]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2044:2040]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2049:2045]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2054:2050]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2069:2065]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2074:2070]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_394_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_394_nl = nl_ACCUM_INNER_LOOP_acc_394_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2079:2075]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2084:2080]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2089:2085]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2094:2090]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_390_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_390_nl = nl_ACCUM_INNER_LOOP_acc_390_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1698_nl = (ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[149:145]);
  assign ACCUM_INNER_LOOP_acc_1698_nl = nl_ACCUM_INNER_LOOP_acc_1698_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2034:2030]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_389_nl = ({ACCUM_INNER_LOOP_acc_1698_nl , (ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_389_nl = nl_ACCUM_INNER_LOOP_acc_389_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_393_nl = ACCUM_INNER_LOOP_acc_390_nl + ACCUM_INNER_LOOP_acc_389_nl;
  assign ACCUM_INNER_LOOP_acc_393_nl = nl_ACCUM_INNER_LOOP_acc_393_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_394_nl
      + ACCUM_INNER_LOOP_acc_393_nl;
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 = (ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2129:2125]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2134:2130]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2109:2105]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2114:2110]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2119:2115]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2124:2120]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2139:2135]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2144:2140]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_407_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_407_nl = nl_ACCUM_INNER_LOOP_acc_407_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2149:2145]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2154:2150]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2159:2155]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2164:2160]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_403_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_403_nl = nl_ACCUM_INNER_LOOP_acc_403_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1699_nl = (ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[154:150]);
  assign ACCUM_INNER_LOOP_acc_1699_nl = nl_ACCUM_INNER_LOOP_acc_1699_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2104:2100]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_402_nl = ({ACCUM_INNER_LOOP_acc_1699_nl , (ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_402_nl = nl_ACCUM_INNER_LOOP_acc_402_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_406_nl = ACCUM_INNER_LOOP_acc_403_nl + ACCUM_INNER_LOOP_acc_402_nl;
  assign ACCUM_INNER_LOOP_acc_406_nl = nl_ACCUM_INNER_LOOP_acc_406_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_407_nl
      + ACCUM_INNER_LOOP_acc_406_nl;
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 = (ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2199:2195]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2204:2200]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2179:2175]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2184:2180]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2189:2185]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2194:2190]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2209:2205]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2214:2210]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_420_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_420_nl = nl_ACCUM_INNER_LOOP_acc_420_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2219:2215]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2224:2220]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2229:2225]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2234:2230]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_416_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_416_nl = nl_ACCUM_INNER_LOOP_acc_416_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1700_nl = (ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[159:155]);
  assign ACCUM_INNER_LOOP_acc_1700_nl = nl_ACCUM_INNER_LOOP_acc_1700_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2174:2170]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_415_nl = ({ACCUM_INNER_LOOP_acc_1700_nl , (ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_415_nl = nl_ACCUM_INNER_LOOP_acc_415_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_419_nl = ACCUM_INNER_LOOP_acc_416_nl + ACCUM_INNER_LOOP_acc_415_nl;
  assign ACCUM_INNER_LOOP_acc_419_nl = nl_ACCUM_INNER_LOOP_acc_419_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_420_nl
      + ACCUM_INNER_LOOP_acc_419_nl;
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 = (ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2269:2265]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2274:2270]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2249:2245]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2254:2250]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2259:2255]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2264:2260]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2279:2275]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2284:2280]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_433_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_433_nl = nl_ACCUM_INNER_LOOP_acc_433_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2289:2285]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2294:2290]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2299:2295]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2304:2300]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_429_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_429_nl = nl_ACCUM_INNER_LOOP_acc_429_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1701_nl = (ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[164:160]);
  assign ACCUM_INNER_LOOP_acc_1701_nl = nl_ACCUM_INNER_LOOP_acc_1701_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2244:2240]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_428_nl = ({ACCUM_INNER_LOOP_acc_1701_nl , (ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_428_nl = nl_ACCUM_INNER_LOOP_acc_428_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_432_nl = ACCUM_INNER_LOOP_acc_429_nl + ACCUM_INNER_LOOP_acc_428_nl;
  assign ACCUM_INNER_LOOP_acc_432_nl = nl_ACCUM_INNER_LOOP_acc_432_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_433_nl
      + ACCUM_INNER_LOOP_acc_432_nl;
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 = (ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2339:2335]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2344:2340]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2319:2315]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2324:2320]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2329:2325]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2334:2330]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2349:2345]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2354:2350]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_446_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_446_nl = nl_ACCUM_INNER_LOOP_acc_446_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2359:2355]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2364:2360]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2369:2365]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2374:2370]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_442_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_442_nl = nl_ACCUM_INNER_LOOP_acc_442_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1702_nl = (ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[169:165]);
  assign ACCUM_INNER_LOOP_acc_1702_nl = nl_ACCUM_INNER_LOOP_acc_1702_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2314:2310]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_441_nl = ({ACCUM_INNER_LOOP_acc_1702_nl , (ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_441_nl = nl_ACCUM_INNER_LOOP_acc_441_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_445_nl = ACCUM_INNER_LOOP_acc_442_nl + ACCUM_INNER_LOOP_acc_441_nl;
  assign ACCUM_INNER_LOOP_acc_445_nl = nl_ACCUM_INNER_LOOP_acc_445_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_446_nl
      + ACCUM_INNER_LOOP_acc_445_nl;
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 = (ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2409:2405]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2414:2410]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2389:2385]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2394:2390]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2399:2395]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2404:2400]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2419:2415]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2424:2420]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_459_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_459_nl = nl_ACCUM_INNER_LOOP_acc_459_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2429:2425]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2434:2430]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2439:2435]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2444:2440]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_455_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_455_nl = nl_ACCUM_INNER_LOOP_acc_455_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1703_nl = (ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[174:170]);
  assign ACCUM_INNER_LOOP_acc_1703_nl = nl_ACCUM_INNER_LOOP_acc_1703_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2384:2380]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_454_nl = ({ACCUM_INNER_LOOP_acc_1703_nl , (ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_454_nl = nl_ACCUM_INNER_LOOP_acc_454_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_458_nl = ACCUM_INNER_LOOP_acc_455_nl + ACCUM_INNER_LOOP_acc_454_nl;
  assign ACCUM_INNER_LOOP_acc_458_nl = nl_ACCUM_INNER_LOOP_acc_458_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_459_nl
      + ACCUM_INNER_LOOP_acc_458_nl;
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 = (ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2479:2475]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2484:2480]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2459:2455]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2464:2460]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2469:2465]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2474:2470]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2489:2485]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2494:2490]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_472_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_472_nl = nl_ACCUM_INNER_LOOP_acc_472_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2499:2495]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2504:2500]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2509:2505]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2514:2510]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_468_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_468_nl = nl_ACCUM_INNER_LOOP_acc_468_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1704_nl = (ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[179:175]);
  assign ACCUM_INNER_LOOP_acc_1704_nl = nl_ACCUM_INNER_LOOP_acc_1704_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2454:2450]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_467_nl = ({ACCUM_INNER_LOOP_acc_1704_nl , (ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_467_nl = nl_ACCUM_INNER_LOOP_acc_467_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_471_nl = ACCUM_INNER_LOOP_acc_468_nl + ACCUM_INNER_LOOP_acc_467_nl;
  assign ACCUM_INNER_LOOP_acc_471_nl = nl_ACCUM_INNER_LOOP_acc_471_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_472_nl
      + ACCUM_INNER_LOOP_acc_471_nl;
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 = (ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2549:2545]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2554:2550]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2529:2525]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2534:2530]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2539:2535]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2544:2540]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2559:2555]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2564:2560]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_485_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_485_nl = nl_ACCUM_INNER_LOOP_acc_485_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2569:2565]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2574:2570]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2579:2575]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2584:2580]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_481_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_481_nl = nl_ACCUM_INNER_LOOP_acc_481_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1705_nl = (ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[184:180]);
  assign ACCUM_INNER_LOOP_acc_1705_nl = nl_ACCUM_INNER_LOOP_acc_1705_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2524:2520]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_480_nl = ({ACCUM_INNER_LOOP_acc_1705_nl , (ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_480_nl = nl_ACCUM_INNER_LOOP_acc_480_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_484_nl = ACCUM_INNER_LOOP_acc_481_nl + ACCUM_INNER_LOOP_acc_480_nl;
  assign ACCUM_INNER_LOOP_acc_484_nl = nl_ACCUM_INNER_LOOP_acc_484_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_485_nl
      + ACCUM_INNER_LOOP_acc_484_nl;
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 = (ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2619:2615]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2624:2620]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2599:2595]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2604:2600]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2609:2605]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2614:2610]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2629:2625]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2634:2630]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_498_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_498_nl = nl_ACCUM_INNER_LOOP_acc_498_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2639:2635]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2644:2640]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2649:2645]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2654:2650]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_494_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_494_nl = nl_ACCUM_INNER_LOOP_acc_494_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1706_nl = (ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[189:185]);
  assign ACCUM_INNER_LOOP_acc_1706_nl = nl_ACCUM_INNER_LOOP_acc_1706_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2594:2590]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_493_nl = ({ACCUM_INNER_LOOP_acc_1706_nl , (ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_493_nl = nl_ACCUM_INNER_LOOP_acc_493_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_497_nl = ACCUM_INNER_LOOP_acc_494_nl + ACCUM_INNER_LOOP_acc_493_nl;
  assign ACCUM_INNER_LOOP_acc_497_nl = nl_ACCUM_INNER_LOOP_acc_497_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_498_nl
      + ACCUM_INNER_LOOP_acc_497_nl;
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 = (ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2689:2685]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2694:2690]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2669:2665]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2674:2670]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2679:2675]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2684:2680]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2699:2695]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2704:2700]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_511_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_511_nl = nl_ACCUM_INNER_LOOP_acc_511_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2709:2705]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2714:2710]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2719:2715]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2724:2720]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_507_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_507_nl = nl_ACCUM_INNER_LOOP_acc_507_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1707_nl = (ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[194:190]);
  assign ACCUM_INNER_LOOP_acc_1707_nl = nl_ACCUM_INNER_LOOP_acc_1707_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2664:2660]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_506_nl = ({ACCUM_INNER_LOOP_acc_1707_nl , (ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_506_nl = nl_ACCUM_INNER_LOOP_acc_506_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_510_nl = ACCUM_INNER_LOOP_acc_507_nl + ACCUM_INNER_LOOP_acc_506_nl;
  assign ACCUM_INNER_LOOP_acc_510_nl = nl_ACCUM_INNER_LOOP_acc_510_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_511_nl
      + ACCUM_INNER_LOOP_acc_510_nl;
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 = (ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2759:2755]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2764:2760]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2739:2735]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2744:2740]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2749:2745]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2754:2750]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2769:2765]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2774:2770]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_524_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_524_nl = nl_ACCUM_INNER_LOOP_acc_524_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2779:2775]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2784:2780]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2789:2785]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2794:2790]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_520_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_520_nl = nl_ACCUM_INNER_LOOP_acc_520_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1708_nl = (ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[199:195]);
  assign ACCUM_INNER_LOOP_acc_1708_nl = nl_ACCUM_INNER_LOOP_acc_1708_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2734:2730]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_519_nl = ({ACCUM_INNER_LOOP_acc_1708_nl , (ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_519_nl = nl_ACCUM_INNER_LOOP_acc_519_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_523_nl = ACCUM_INNER_LOOP_acc_520_nl + ACCUM_INNER_LOOP_acc_519_nl;
  assign ACCUM_INNER_LOOP_acc_523_nl = nl_ACCUM_INNER_LOOP_acc_523_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_524_nl
      + ACCUM_INNER_LOOP_acc_523_nl;
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 = (ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2829:2825]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2834:2830]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2809:2805]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2814:2810]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2819:2815]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2824:2820]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2839:2835]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2844:2840]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_537_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_537_nl = nl_ACCUM_INNER_LOOP_acc_537_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2849:2845]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2854:2850]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2859:2855]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2864:2860]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_533_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_533_nl = nl_ACCUM_INNER_LOOP_acc_533_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1709_nl = (ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[204:200]);
  assign ACCUM_INNER_LOOP_acc_1709_nl = nl_ACCUM_INNER_LOOP_acc_1709_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2804:2800]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_532_nl = ({ACCUM_INNER_LOOP_acc_1709_nl , (ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_532_nl = nl_ACCUM_INNER_LOOP_acc_532_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_536_nl = ACCUM_INNER_LOOP_acc_533_nl + ACCUM_INNER_LOOP_acc_532_nl;
  assign ACCUM_INNER_LOOP_acc_536_nl = nl_ACCUM_INNER_LOOP_acc_536_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_537_nl
      + ACCUM_INNER_LOOP_acc_536_nl;
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 = (ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2899:2895]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2904:2900]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2879:2875]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2884:2880]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2889:2885]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2894:2890]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2909:2905]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2914:2910]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_550_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_550_nl = nl_ACCUM_INNER_LOOP_acc_550_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2919:2915]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2924:2920]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2929:2925]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[2934:2930]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_546_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_546_nl = nl_ACCUM_INNER_LOOP_acc_546_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1710_nl = (ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[209:205]);
  assign ACCUM_INNER_LOOP_acc_1710_nl = nl_ACCUM_INNER_LOOP_acc_1710_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2874:2870]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_545_nl = ({ACCUM_INNER_LOOP_acc_1710_nl , (ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_545_nl = nl_ACCUM_INNER_LOOP_acc_545_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_549_nl = ACCUM_INNER_LOOP_acc_546_nl + ACCUM_INNER_LOOP_acc_545_nl;
  assign ACCUM_INNER_LOOP_acc_549_nl = nl_ACCUM_INNER_LOOP_acc_549_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_550_nl
      + ACCUM_INNER_LOOP_acc_549_nl;
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 = (ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[2969:2965]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[2974:2970]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[2949:2945]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[2954:2950]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[2959:2955]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[2964:2960]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[2979:2975]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[2984:2980]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_563_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_563_nl = nl_ACCUM_INNER_LOOP_acc_563_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[2989:2985]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[2994:2990]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[2999:2995]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3004:3000]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_559_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_559_nl = nl_ACCUM_INNER_LOOP_acc_559_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1711_nl = (ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[214:210]);
  assign ACCUM_INNER_LOOP_acc_1711_nl = nl_ACCUM_INNER_LOOP_acc_1711_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[2944:2940]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_558_nl = ({ACCUM_INNER_LOOP_acc_1711_nl , (ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_558_nl = nl_ACCUM_INNER_LOOP_acc_558_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_562_nl = ACCUM_INNER_LOOP_acc_559_nl + ACCUM_INNER_LOOP_acc_558_nl;
  assign ACCUM_INNER_LOOP_acc_562_nl = nl_ACCUM_INNER_LOOP_acc_562_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_563_nl
      + ACCUM_INNER_LOOP_acc_562_nl;
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 = (ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3039:3035]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3044:3040]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3019:3015]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3024:3020]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3029:3025]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3034:3030]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3049:3045]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3054:3050]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_576_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_576_nl = nl_ACCUM_INNER_LOOP_acc_576_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3059:3055]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3064:3060]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3069:3065]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3074:3070]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_572_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_572_nl = nl_ACCUM_INNER_LOOP_acc_572_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1712_nl = (ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[219:215]);
  assign ACCUM_INNER_LOOP_acc_1712_nl = nl_ACCUM_INNER_LOOP_acc_1712_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3014:3010]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_571_nl = ({ACCUM_INNER_LOOP_acc_1712_nl , (ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_571_nl = nl_ACCUM_INNER_LOOP_acc_571_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_575_nl = ACCUM_INNER_LOOP_acc_572_nl + ACCUM_INNER_LOOP_acc_571_nl;
  assign ACCUM_INNER_LOOP_acc_575_nl = nl_ACCUM_INNER_LOOP_acc_575_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_576_nl
      + ACCUM_INNER_LOOP_acc_575_nl;
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 = (ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3109:3105]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3114:3110]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3089:3085]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3094:3090]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3099:3095]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3104:3100]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3119:3115]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3124:3120]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_589_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_589_nl = nl_ACCUM_INNER_LOOP_acc_589_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3129:3125]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3134:3130]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3139:3135]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3144:3140]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_585_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_585_nl = nl_ACCUM_INNER_LOOP_acc_585_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1713_nl = (ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[224:220]);
  assign ACCUM_INNER_LOOP_acc_1713_nl = nl_ACCUM_INNER_LOOP_acc_1713_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3084:3080]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_584_nl = ({ACCUM_INNER_LOOP_acc_1713_nl , (ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_584_nl = nl_ACCUM_INNER_LOOP_acc_584_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_588_nl = ACCUM_INNER_LOOP_acc_585_nl + ACCUM_INNER_LOOP_acc_584_nl;
  assign ACCUM_INNER_LOOP_acc_588_nl = nl_ACCUM_INNER_LOOP_acc_588_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_589_nl
      + ACCUM_INNER_LOOP_acc_588_nl;
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 = (ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3179:3175]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3184:3180]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3159:3155]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3164:3160]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3169:3165]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3174:3170]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3189:3185]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3194:3190]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_602_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_602_nl = nl_ACCUM_INNER_LOOP_acc_602_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3199:3195]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3204:3200]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3209:3205]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3214:3210]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_598_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_598_nl = nl_ACCUM_INNER_LOOP_acc_598_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1714_nl = (ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[229:225]);
  assign ACCUM_INNER_LOOP_acc_1714_nl = nl_ACCUM_INNER_LOOP_acc_1714_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3154:3150]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_597_nl = ({ACCUM_INNER_LOOP_acc_1714_nl , (ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_597_nl = nl_ACCUM_INNER_LOOP_acc_597_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_601_nl = ACCUM_INNER_LOOP_acc_598_nl + ACCUM_INNER_LOOP_acc_597_nl;
  assign ACCUM_INNER_LOOP_acc_601_nl = nl_ACCUM_INNER_LOOP_acc_601_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_602_nl
      + ACCUM_INNER_LOOP_acc_601_nl;
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 = (ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3249:3245]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3254:3250]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3229:3225]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3234:3230]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3239:3235]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3244:3240]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3259:3255]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3264:3260]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_615_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_615_nl = nl_ACCUM_INNER_LOOP_acc_615_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3269:3265]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3274:3270]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3279:3275]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3284:3280]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_611_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_611_nl = nl_ACCUM_INNER_LOOP_acc_611_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1715_nl = (ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[234:230]);
  assign ACCUM_INNER_LOOP_acc_1715_nl = nl_ACCUM_INNER_LOOP_acc_1715_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3224:3220]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_610_nl = ({ACCUM_INNER_LOOP_acc_1715_nl , (ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_610_nl = nl_ACCUM_INNER_LOOP_acc_610_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_614_nl = ACCUM_INNER_LOOP_acc_611_nl + ACCUM_INNER_LOOP_acc_610_nl;
  assign ACCUM_INNER_LOOP_acc_614_nl = nl_ACCUM_INNER_LOOP_acc_614_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_615_nl
      + ACCUM_INNER_LOOP_acc_614_nl;
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 = (ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3319:3315]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3324:3320]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3299:3295]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3304:3300]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3309:3305]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3314:3310]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3329:3325]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3334:3330]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_628_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_628_nl = nl_ACCUM_INNER_LOOP_acc_628_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3339:3335]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3344:3340]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3349:3345]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3354:3350]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_624_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_624_nl = nl_ACCUM_INNER_LOOP_acc_624_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1716_nl = (ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[239:235]);
  assign ACCUM_INNER_LOOP_acc_1716_nl = nl_ACCUM_INNER_LOOP_acc_1716_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3294:3290]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_623_nl = ({ACCUM_INNER_LOOP_acc_1716_nl , (ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_623_nl = nl_ACCUM_INNER_LOOP_acc_623_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_627_nl = ACCUM_INNER_LOOP_acc_624_nl + ACCUM_INNER_LOOP_acc_623_nl;
  assign ACCUM_INNER_LOOP_acc_627_nl = nl_ACCUM_INNER_LOOP_acc_627_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_628_nl
      + ACCUM_INNER_LOOP_acc_627_nl;
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 = (ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3389:3385]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3394:3390]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3369:3365]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3374:3370]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3379:3375]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3384:3380]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3399:3395]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3404:3400]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_641_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_641_nl = nl_ACCUM_INNER_LOOP_acc_641_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3409:3405]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3414:3410]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3419:3415]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3424:3420]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_637_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_637_nl = nl_ACCUM_INNER_LOOP_acc_637_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1717_nl = (ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[244:240]);
  assign ACCUM_INNER_LOOP_acc_1717_nl = nl_ACCUM_INNER_LOOP_acc_1717_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3364:3360]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_636_nl = ({ACCUM_INNER_LOOP_acc_1717_nl , (ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_636_nl = nl_ACCUM_INNER_LOOP_acc_636_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_640_nl = ACCUM_INNER_LOOP_acc_637_nl + ACCUM_INNER_LOOP_acc_636_nl;
  assign ACCUM_INNER_LOOP_acc_640_nl = nl_ACCUM_INNER_LOOP_acc_640_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_641_nl
      + ACCUM_INNER_LOOP_acc_640_nl;
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 = (ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3459:3455]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3464:3460]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3439:3435]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3444:3440]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3449:3445]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3454:3450]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3469:3465]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3474:3470]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_654_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_654_nl = nl_ACCUM_INNER_LOOP_acc_654_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3479:3475]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3484:3480]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3489:3485]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3494:3490]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_650_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_650_nl = nl_ACCUM_INNER_LOOP_acc_650_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1718_nl = (ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[249:245]);
  assign ACCUM_INNER_LOOP_acc_1718_nl = nl_ACCUM_INNER_LOOP_acc_1718_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3434:3430]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_649_nl = ({ACCUM_INNER_LOOP_acc_1718_nl , (ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_649_nl = nl_ACCUM_INNER_LOOP_acc_649_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_653_nl = ACCUM_INNER_LOOP_acc_650_nl + ACCUM_INNER_LOOP_acc_649_nl;
  assign ACCUM_INNER_LOOP_acc_653_nl = nl_ACCUM_INNER_LOOP_acc_653_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_654_nl
      + ACCUM_INNER_LOOP_acc_653_nl;
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 = (ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3529:3525]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3534:3530]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3509:3505]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3514:3510]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3519:3515]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3524:3520]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3539:3535]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3544:3540]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_667_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_667_nl = nl_ACCUM_INNER_LOOP_acc_667_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3549:3545]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3554:3550]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3559:3555]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3564:3560]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_663_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_663_nl = nl_ACCUM_INNER_LOOP_acc_663_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1719_nl = (ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[254:250]);
  assign ACCUM_INNER_LOOP_acc_1719_nl = nl_ACCUM_INNER_LOOP_acc_1719_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3504:3500]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_662_nl = ({ACCUM_INNER_LOOP_acc_1719_nl , (ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_662_nl = nl_ACCUM_INNER_LOOP_acc_662_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_666_nl = ACCUM_INNER_LOOP_acc_663_nl + ACCUM_INNER_LOOP_acc_662_nl;
  assign ACCUM_INNER_LOOP_acc_666_nl = nl_ACCUM_INNER_LOOP_acc_666_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_667_nl
      + ACCUM_INNER_LOOP_acc_666_nl;
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 = (ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3599:3595]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3604:3600]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3579:3575]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3584:3580]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3589:3585]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3594:3590]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3609:3605]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3614:3610]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_680_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_680_nl = nl_ACCUM_INNER_LOOP_acc_680_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3619:3615]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3624:3620]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3629:3625]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3634:3630]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_676_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_676_nl = nl_ACCUM_INNER_LOOP_acc_676_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1720_nl = (ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[259:255]);
  assign ACCUM_INNER_LOOP_acc_1720_nl = nl_ACCUM_INNER_LOOP_acc_1720_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3574:3570]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_675_nl = ({ACCUM_INNER_LOOP_acc_1720_nl , (ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_675_nl = nl_ACCUM_INNER_LOOP_acc_675_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_679_nl = ACCUM_INNER_LOOP_acc_676_nl + ACCUM_INNER_LOOP_acc_675_nl;
  assign ACCUM_INNER_LOOP_acc_679_nl = nl_ACCUM_INNER_LOOP_acc_679_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_680_nl
      + ACCUM_INNER_LOOP_acc_679_nl;
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 = (ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3669:3665]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3674:3670]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3649:3645]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3654:3650]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3659:3655]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3664:3660]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3679:3675]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3684:3680]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_693_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_693_nl = nl_ACCUM_INNER_LOOP_acc_693_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3689:3685]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3694:3690]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3699:3695]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3704:3700]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_689_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_689_nl = nl_ACCUM_INNER_LOOP_acc_689_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1721_nl = (ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[264:260]);
  assign ACCUM_INNER_LOOP_acc_1721_nl = nl_ACCUM_INNER_LOOP_acc_1721_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3644:3640]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_688_nl = ({ACCUM_INNER_LOOP_acc_1721_nl , (ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_688_nl = nl_ACCUM_INNER_LOOP_acc_688_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_692_nl = ACCUM_INNER_LOOP_acc_689_nl + ACCUM_INNER_LOOP_acc_688_nl;
  assign ACCUM_INNER_LOOP_acc_692_nl = nl_ACCUM_INNER_LOOP_acc_692_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_693_nl
      + ACCUM_INNER_LOOP_acc_692_nl;
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 = (ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3739:3735]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3744:3740]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3719:3715]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3724:3720]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3729:3725]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3734:3730]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3749:3745]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3754:3750]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_706_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_706_nl = nl_ACCUM_INNER_LOOP_acc_706_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3759:3755]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3764:3760]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3769:3765]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3774:3770]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_702_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_702_nl = nl_ACCUM_INNER_LOOP_acc_702_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1722_nl = (ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[269:265]);
  assign ACCUM_INNER_LOOP_acc_1722_nl = nl_ACCUM_INNER_LOOP_acc_1722_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3714:3710]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_701_nl = ({ACCUM_INNER_LOOP_acc_1722_nl , (ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_701_nl = nl_ACCUM_INNER_LOOP_acc_701_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_705_nl = ACCUM_INNER_LOOP_acc_702_nl + ACCUM_INNER_LOOP_acc_701_nl;
  assign ACCUM_INNER_LOOP_acc_705_nl = nl_ACCUM_INNER_LOOP_acc_705_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_706_nl
      + ACCUM_INNER_LOOP_acc_705_nl;
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 = (ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3809:3805]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3814:3810]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3789:3785]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3794:3790]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3799:3795]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3804:3800]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3819:3815]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3824:3820]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_719_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_719_nl = nl_ACCUM_INNER_LOOP_acc_719_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3829:3825]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3834:3830]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3839:3835]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3844:3840]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_715_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_715_nl = nl_ACCUM_INNER_LOOP_acc_715_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1723_nl = (ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[274:270]);
  assign ACCUM_INNER_LOOP_acc_1723_nl = nl_ACCUM_INNER_LOOP_acc_1723_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3784:3780]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_714_nl = ({ACCUM_INNER_LOOP_acc_1723_nl , (ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_714_nl = nl_ACCUM_INNER_LOOP_acc_714_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_718_nl = ACCUM_INNER_LOOP_acc_715_nl + ACCUM_INNER_LOOP_acc_714_nl;
  assign ACCUM_INNER_LOOP_acc_718_nl = nl_ACCUM_INNER_LOOP_acc_718_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_719_nl
      + ACCUM_INNER_LOOP_acc_718_nl;
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 = (ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3879:3875]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3884:3880]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3859:3855]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3864:3860]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3869:3865]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3874:3870]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3889:3885]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3894:3890]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_732_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_732_nl = nl_ACCUM_INNER_LOOP_acc_732_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3899:3895]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3904:3900]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3909:3905]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3914:3910]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_728_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_728_nl = nl_ACCUM_INNER_LOOP_acc_728_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1724_nl = (ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[279:275]);
  assign ACCUM_INNER_LOOP_acc_1724_nl = nl_ACCUM_INNER_LOOP_acc_1724_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3854:3850]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_727_nl = ({ACCUM_INNER_LOOP_acc_1724_nl , (ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_727_nl = nl_ACCUM_INNER_LOOP_acc_727_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_731_nl = ACCUM_INNER_LOOP_acc_728_nl + ACCUM_INNER_LOOP_acc_727_nl;
  assign ACCUM_INNER_LOOP_acc_731_nl = nl_ACCUM_INNER_LOOP_acc_731_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_732_nl
      + ACCUM_INNER_LOOP_acc_731_nl;
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 = (ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[3949:3945]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[3954:3950]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3929:3925]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[3934:3930]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[3939:3935]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[3944:3940]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[3959:3955]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[3964:3960]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_745_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_745_nl = nl_ACCUM_INNER_LOOP_acc_745_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[3969:3965]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[3974:3970]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[3979:3975]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[3984:3980]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_741_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_741_nl = nl_ACCUM_INNER_LOOP_acc_741_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1725_nl = (ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[284:280]);
  assign ACCUM_INNER_LOOP_acc_1725_nl = nl_ACCUM_INNER_LOOP_acc_1725_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3924:3920]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_740_nl = ({ACCUM_INNER_LOOP_acc_1725_nl , (ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_740_nl = nl_ACCUM_INNER_LOOP_acc_740_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_744_nl = ACCUM_INNER_LOOP_acc_741_nl + ACCUM_INNER_LOOP_acc_740_nl;
  assign ACCUM_INNER_LOOP_acc_744_nl = nl_ACCUM_INNER_LOOP_acc_744_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_745_nl
      + ACCUM_INNER_LOOP_acc_744_nl;
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1 = (ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4019:4015]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4024:4020]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[3999:3995]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4004:4000]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4009:4005]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4014:4010]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4029:4025]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4034:4030]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_758_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_758_nl = nl_ACCUM_INNER_LOOP_acc_758_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4039:4035]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4044:4040]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4049:4045]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4054:4050]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_754_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_754_nl = nl_ACCUM_INNER_LOOP_acc_754_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1726_nl = (ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[289:285]);
  assign ACCUM_INNER_LOOP_acc_1726_nl = nl_ACCUM_INNER_LOOP_acc_1726_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[3994:3990]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_753_nl = ({ACCUM_INNER_LOOP_acc_1726_nl , (ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_753_nl = nl_ACCUM_INNER_LOOP_acc_753_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_757_nl = ACCUM_INNER_LOOP_acc_754_nl + ACCUM_INNER_LOOP_acc_753_nl;
  assign ACCUM_INNER_LOOP_acc_757_nl = nl_ACCUM_INNER_LOOP_acc_757_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_758_nl
      + ACCUM_INNER_LOOP_acc_757_nl;
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1 = (ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4089:4085]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4094:4090]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4069:4065]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4074:4070]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4079:4075]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4084:4080]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4099:4095]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4104:4100]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_771_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_771_nl = nl_ACCUM_INNER_LOOP_acc_771_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4109:4105]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4114:4110]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4119:4115]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4124:4120]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_767_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_767_nl = nl_ACCUM_INNER_LOOP_acc_767_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1727_nl = (ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[294:290]);
  assign ACCUM_INNER_LOOP_acc_1727_nl = nl_ACCUM_INNER_LOOP_acc_1727_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4064:4060]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_766_nl = ({ACCUM_INNER_LOOP_acc_1727_nl , (ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_766_nl = nl_ACCUM_INNER_LOOP_acc_766_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_770_nl = ACCUM_INNER_LOOP_acc_767_nl + ACCUM_INNER_LOOP_acc_766_nl;
  assign ACCUM_INNER_LOOP_acc_770_nl = nl_ACCUM_INNER_LOOP_acc_770_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_771_nl
      + ACCUM_INNER_LOOP_acc_770_nl;
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1 = (ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4159:4155]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4164:4160]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4139:4135]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4144:4140]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4149:4145]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4154:4150]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4169:4165]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4174:4170]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_784_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_784_nl = nl_ACCUM_INNER_LOOP_acc_784_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4179:4175]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4184:4180]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4189:4185]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4194:4190]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_780_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_780_nl = nl_ACCUM_INNER_LOOP_acc_780_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1728_nl = (ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[299:295]);
  assign ACCUM_INNER_LOOP_acc_1728_nl = nl_ACCUM_INNER_LOOP_acc_1728_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4134:4130]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_779_nl = ({ACCUM_INNER_LOOP_acc_1728_nl , (ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_779_nl = nl_ACCUM_INNER_LOOP_acc_779_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_783_nl = ACCUM_INNER_LOOP_acc_780_nl + ACCUM_INNER_LOOP_acc_779_nl;
  assign ACCUM_INNER_LOOP_acc_783_nl = nl_ACCUM_INNER_LOOP_acc_783_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_784_nl
      + ACCUM_INNER_LOOP_acc_783_nl;
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1 = (ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4229:4225]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4234:4230]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4209:4205]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4214:4210]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4219:4215]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4224:4220]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4239:4235]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4244:4240]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_797_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_797_nl = nl_ACCUM_INNER_LOOP_acc_797_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4249:4245]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4254:4250]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4259:4255]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4264:4260]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_793_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_793_nl = nl_ACCUM_INNER_LOOP_acc_793_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1729_nl = (ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[304:300]);
  assign ACCUM_INNER_LOOP_acc_1729_nl = nl_ACCUM_INNER_LOOP_acc_1729_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4204:4200]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_792_nl = ({ACCUM_INNER_LOOP_acc_1729_nl , (ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_792_nl = nl_ACCUM_INNER_LOOP_acc_792_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_796_nl = ACCUM_INNER_LOOP_acc_793_nl + ACCUM_INNER_LOOP_acc_792_nl;
  assign ACCUM_INNER_LOOP_acc_796_nl = nl_ACCUM_INNER_LOOP_acc_796_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_797_nl
      + ACCUM_INNER_LOOP_acc_796_nl;
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1 = (ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4299:4295]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4304:4300]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4279:4275]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4284:4280]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4289:4285]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4294:4290]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4309:4305]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4314:4310]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_810_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_810_nl = nl_ACCUM_INNER_LOOP_acc_810_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4319:4315]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4324:4320]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4329:4325]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4334:4330]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_806_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_806_nl = nl_ACCUM_INNER_LOOP_acc_806_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1730_nl = (ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[309:305]);
  assign ACCUM_INNER_LOOP_acc_1730_nl = nl_ACCUM_INNER_LOOP_acc_1730_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4274:4270]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_805_nl = ({ACCUM_INNER_LOOP_acc_1730_nl , (ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_805_nl = nl_ACCUM_INNER_LOOP_acc_805_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_809_nl = ACCUM_INNER_LOOP_acc_806_nl + ACCUM_INNER_LOOP_acc_805_nl;
  assign ACCUM_INNER_LOOP_acc_809_nl = nl_ACCUM_INNER_LOOP_acc_809_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_810_nl
      + ACCUM_INNER_LOOP_acc_809_nl;
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1 = (ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4369:4365]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4374:4370]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4349:4345]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4354:4350]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4359:4355]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4364:4360]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4379:4375]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4384:4380]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_823_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_823_nl = nl_ACCUM_INNER_LOOP_acc_823_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4389:4385]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4394:4390]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4399:4395]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4404:4400]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_819_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_819_nl = nl_ACCUM_INNER_LOOP_acc_819_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1731_nl = (ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[314:310]);
  assign ACCUM_INNER_LOOP_acc_1731_nl = nl_ACCUM_INNER_LOOP_acc_1731_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4344:4340]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_818_nl = ({ACCUM_INNER_LOOP_acc_1731_nl , (ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_818_nl = nl_ACCUM_INNER_LOOP_acc_818_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_822_nl = ACCUM_INNER_LOOP_acc_819_nl + ACCUM_INNER_LOOP_acc_818_nl;
  assign ACCUM_INNER_LOOP_acc_822_nl = nl_ACCUM_INNER_LOOP_acc_822_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_823_nl
      + ACCUM_INNER_LOOP_acc_822_nl;
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1 = (ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4439:4435]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4444:4440]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4419:4415]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4424:4420]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4429:4425]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4434:4430]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4449:4445]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4454:4450]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_836_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_836_nl = nl_ACCUM_INNER_LOOP_acc_836_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4459:4455]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4464:4460]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4469:4465]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4474:4470]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_832_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_832_nl = nl_ACCUM_INNER_LOOP_acc_832_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1732_nl = (ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[319:315]);
  assign ACCUM_INNER_LOOP_acc_1732_nl = nl_ACCUM_INNER_LOOP_acc_1732_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4414:4410]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_831_nl = ({ACCUM_INNER_LOOP_acc_1732_nl , (ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_831_nl = nl_ACCUM_INNER_LOOP_acc_831_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_835_nl = ACCUM_INNER_LOOP_acc_832_nl + ACCUM_INNER_LOOP_acc_831_nl;
  assign ACCUM_INNER_LOOP_acc_835_nl = nl_ACCUM_INNER_LOOP_acc_835_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_836_nl
      + ACCUM_INNER_LOOP_acc_835_nl;
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1 = (ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4509:4505]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4514:4510]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4489:4485]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4494:4490]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4499:4495]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4504:4500]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4519:4515]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4524:4520]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_849_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_849_nl = nl_ACCUM_INNER_LOOP_acc_849_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4529:4525]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4534:4530]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4539:4535]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4544:4540]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_845_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_845_nl = nl_ACCUM_INNER_LOOP_acc_845_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1733_nl = (ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[324:320]);
  assign ACCUM_INNER_LOOP_acc_1733_nl = nl_ACCUM_INNER_LOOP_acc_1733_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4484:4480]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_844_nl = ({ACCUM_INNER_LOOP_acc_1733_nl , (ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_844_nl = nl_ACCUM_INNER_LOOP_acc_844_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_848_nl = ACCUM_INNER_LOOP_acc_845_nl + ACCUM_INNER_LOOP_acc_844_nl;
  assign ACCUM_INNER_LOOP_acc_848_nl = nl_ACCUM_INNER_LOOP_acc_848_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_849_nl
      + ACCUM_INNER_LOOP_acc_848_nl;
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1 = (ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4579:4575]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4584:4580]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4559:4555]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4564:4560]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4569:4565]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4574:4570]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4589:4585]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4594:4590]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_862_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_862_nl = nl_ACCUM_INNER_LOOP_acc_862_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4599:4595]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4604:4600]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4609:4605]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4614:4610]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_858_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_858_nl = nl_ACCUM_INNER_LOOP_acc_858_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1734_nl = (ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[329:325]);
  assign ACCUM_INNER_LOOP_acc_1734_nl = nl_ACCUM_INNER_LOOP_acc_1734_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4554:4550]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_857_nl = ({ACCUM_INNER_LOOP_acc_1734_nl , (ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_857_nl = nl_ACCUM_INNER_LOOP_acc_857_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_861_nl = ACCUM_INNER_LOOP_acc_858_nl + ACCUM_INNER_LOOP_acc_857_nl;
  assign ACCUM_INNER_LOOP_acc_861_nl = nl_ACCUM_INNER_LOOP_acc_861_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_862_nl
      + ACCUM_INNER_LOOP_acc_861_nl;
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1 = (ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4649:4645]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4654:4650]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4629:4625]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4634:4630]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4639:4635]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4644:4640]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4659:4655]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4664:4660]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_875_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_875_nl = nl_ACCUM_INNER_LOOP_acc_875_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4669:4665]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4674:4670]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4679:4675]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4684:4680]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_871_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_871_nl = nl_ACCUM_INNER_LOOP_acc_871_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1735_nl = (ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[334:330]);
  assign ACCUM_INNER_LOOP_acc_1735_nl = nl_ACCUM_INNER_LOOP_acc_1735_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4624:4620]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_870_nl = ({ACCUM_INNER_LOOP_acc_1735_nl , (ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_870_nl = nl_ACCUM_INNER_LOOP_acc_870_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_874_nl = ACCUM_INNER_LOOP_acc_871_nl + ACCUM_INNER_LOOP_acc_870_nl;
  assign ACCUM_INNER_LOOP_acc_874_nl = nl_ACCUM_INNER_LOOP_acc_874_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_875_nl
      + ACCUM_INNER_LOOP_acc_874_nl;
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1 = (ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4719:4715]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4724:4720]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4699:4695]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4704:4700]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4709:4705]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4714:4710]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4729:4725]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4734:4730]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_888_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_888_nl = nl_ACCUM_INNER_LOOP_acc_888_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4739:4735]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4744:4740]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4749:4745]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4754:4750]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_884_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_884_nl = nl_ACCUM_INNER_LOOP_acc_884_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1736_nl = (ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[339:335]);
  assign ACCUM_INNER_LOOP_acc_1736_nl = nl_ACCUM_INNER_LOOP_acc_1736_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4694:4690]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_883_nl = ({ACCUM_INNER_LOOP_acc_1736_nl , (ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_883_nl = nl_ACCUM_INNER_LOOP_acc_883_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_887_nl = ACCUM_INNER_LOOP_acc_884_nl + ACCUM_INNER_LOOP_acc_883_nl;
  assign ACCUM_INNER_LOOP_acc_887_nl = nl_ACCUM_INNER_LOOP_acc_887_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_888_nl
      + ACCUM_INNER_LOOP_acc_887_nl;
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1 = (ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4789:4785]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4794:4790]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4769:4765]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4774:4770]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4779:4775]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4784:4780]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4799:4795]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4804:4800]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_901_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_901_nl = nl_ACCUM_INNER_LOOP_acc_901_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4809:4805]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4814:4810]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4819:4815]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4824:4820]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_897_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_897_nl = nl_ACCUM_INNER_LOOP_acc_897_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1737_nl = (ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[344:340]);
  assign ACCUM_INNER_LOOP_acc_1737_nl = nl_ACCUM_INNER_LOOP_acc_1737_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4764:4760]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_896_nl = ({ACCUM_INNER_LOOP_acc_1737_nl , (ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_896_nl = nl_ACCUM_INNER_LOOP_acc_896_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_900_nl = ACCUM_INNER_LOOP_acc_897_nl + ACCUM_INNER_LOOP_acc_896_nl;
  assign ACCUM_INNER_LOOP_acc_900_nl = nl_ACCUM_INNER_LOOP_acc_900_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_901_nl
      + ACCUM_INNER_LOOP_acc_900_nl;
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1 = (ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4859:4855]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4864:4860]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4839:4835]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4844:4840]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4849:4845]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4854:4850]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4869:4865]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4874:4870]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_914_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_914_nl = nl_ACCUM_INNER_LOOP_acc_914_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4879:4875]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4884:4880]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4889:4885]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4894:4890]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_910_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_910_nl = nl_ACCUM_INNER_LOOP_acc_910_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1738_nl = (ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[349:345]);
  assign ACCUM_INNER_LOOP_acc_1738_nl = nl_ACCUM_INNER_LOOP_acc_1738_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4834:4830]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_909_nl = ({ACCUM_INNER_LOOP_acc_1738_nl , (ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_909_nl = nl_ACCUM_INNER_LOOP_acc_909_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_913_nl = ACCUM_INNER_LOOP_acc_910_nl + ACCUM_INNER_LOOP_acc_909_nl;
  assign ACCUM_INNER_LOOP_acc_913_nl = nl_ACCUM_INNER_LOOP_acc_913_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_914_nl
      + ACCUM_INNER_LOOP_acc_913_nl;
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1 = (ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4929:4925]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[4934:4930]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4909:4905]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4914:4910]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4919:4915]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4924:4920]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[4939:4935]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[4944:4940]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_927_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_927_nl = nl_ACCUM_INNER_LOOP_acc_927_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[4949:4945]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[4954:4950]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[4959:4955]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[4964:4960]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_923_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_923_nl = nl_ACCUM_INNER_LOOP_acc_923_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1739_nl = (ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[354:350]);
  assign ACCUM_INNER_LOOP_acc_1739_nl = nl_ACCUM_INNER_LOOP_acc_1739_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4904:4900]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_922_nl = ({ACCUM_INNER_LOOP_acc_1739_nl , (ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_922_nl = nl_ACCUM_INNER_LOOP_acc_922_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_926_nl = ACCUM_INNER_LOOP_acc_923_nl + ACCUM_INNER_LOOP_acc_922_nl;
  assign ACCUM_INNER_LOOP_acc_926_nl = nl_ACCUM_INNER_LOOP_acc_926_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_927_nl
      + ACCUM_INNER_LOOP_acc_926_nl;
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1 = (ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[4999:4995]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5004:5000]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[4979:4975]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[4984:4980]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[4989:4985]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[4994:4990]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5009:5005]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5014:5010]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_940_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_940_nl = nl_ACCUM_INNER_LOOP_acc_940_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5019:5015]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5024:5020]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5029:5025]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5034:5030]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_936_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_936_nl = nl_ACCUM_INNER_LOOP_acc_936_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1740_nl = (ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[359:355]);
  assign ACCUM_INNER_LOOP_acc_1740_nl = nl_ACCUM_INNER_LOOP_acc_1740_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[4974:4970]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_935_nl = ({ACCUM_INNER_LOOP_acc_1740_nl , (ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_935_nl = nl_ACCUM_INNER_LOOP_acc_935_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_939_nl = ACCUM_INNER_LOOP_acc_936_nl + ACCUM_INNER_LOOP_acc_935_nl;
  assign ACCUM_INNER_LOOP_acc_939_nl = nl_ACCUM_INNER_LOOP_acc_939_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_940_nl
      + ACCUM_INNER_LOOP_acc_939_nl;
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1 = (ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5069:5065]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5074:5070]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5049:5045]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5054:5050]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5059:5055]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5064:5060]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5079:5075]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5084:5080]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_953_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_953_nl = nl_ACCUM_INNER_LOOP_acc_953_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5089:5085]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5094:5090]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5099:5095]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5104:5100]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_949_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_949_nl = nl_ACCUM_INNER_LOOP_acc_949_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1741_nl = (ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[364:360]);
  assign ACCUM_INNER_LOOP_acc_1741_nl = nl_ACCUM_INNER_LOOP_acc_1741_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5044:5040]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_948_nl = ({ACCUM_INNER_LOOP_acc_1741_nl , (ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_948_nl = nl_ACCUM_INNER_LOOP_acc_948_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_952_nl = ACCUM_INNER_LOOP_acc_949_nl + ACCUM_INNER_LOOP_acc_948_nl;
  assign ACCUM_INNER_LOOP_acc_952_nl = nl_ACCUM_INNER_LOOP_acc_952_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_953_nl
      + ACCUM_INNER_LOOP_acc_952_nl;
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1 = (ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5139:5135]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5144:5140]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5119:5115]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5124:5120]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5129:5125]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5134:5130]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5149:5145]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5154:5150]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_966_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_966_nl = nl_ACCUM_INNER_LOOP_acc_966_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5159:5155]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5164:5160]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5169:5165]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5174:5170]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_962_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_962_nl = nl_ACCUM_INNER_LOOP_acc_962_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1742_nl = (ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[369:365]);
  assign ACCUM_INNER_LOOP_acc_1742_nl = nl_ACCUM_INNER_LOOP_acc_1742_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5114:5110]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_961_nl = ({ACCUM_INNER_LOOP_acc_1742_nl , (ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_961_nl = nl_ACCUM_INNER_LOOP_acc_961_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_965_nl = ACCUM_INNER_LOOP_acc_962_nl + ACCUM_INNER_LOOP_acc_961_nl;
  assign ACCUM_INNER_LOOP_acc_965_nl = nl_ACCUM_INNER_LOOP_acc_965_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_966_nl
      + ACCUM_INNER_LOOP_acc_965_nl;
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1 = (ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5209:5205]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5214:5210]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5189:5185]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5194:5190]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5199:5195]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5204:5200]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5219:5215]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5224:5220]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_979_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_979_nl = nl_ACCUM_INNER_LOOP_acc_979_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5229:5225]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5234:5230]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5239:5235]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5244:5240]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_975_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_975_nl = nl_ACCUM_INNER_LOOP_acc_975_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1743_nl = (ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[374:370]);
  assign ACCUM_INNER_LOOP_acc_1743_nl = nl_ACCUM_INNER_LOOP_acc_1743_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5184:5180]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_974_nl = ({ACCUM_INNER_LOOP_acc_1743_nl , (ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_974_nl = nl_ACCUM_INNER_LOOP_acc_974_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_978_nl = ACCUM_INNER_LOOP_acc_975_nl + ACCUM_INNER_LOOP_acc_974_nl;
  assign ACCUM_INNER_LOOP_acc_978_nl = nl_ACCUM_INNER_LOOP_acc_978_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_979_nl
      + ACCUM_INNER_LOOP_acc_978_nl;
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1 = (ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5279:5275]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5284:5280]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5259:5255]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5264:5260]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5269:5265]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5274:5270]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5289:5285]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5294:5290]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_992_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_992_nl = nl_ACCUM_INNER_LOOP_acc_992_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5299:5295]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5304:5300]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5309:5305]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5314:5310]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_988_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_988_nl = nl_ACCUM_INNER_LOOP_acc_988_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1744_nl = (ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[379:375]);
  assign ACCUM_INNER_LOOP_acc_1744_nl = nl_ACCUM_INNER_LOOP_acc_1744_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5254:5250]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_987_nl = ({ACCUM_INNER_LOOP_acc_1744_nl , (ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_987_nl = nl_ACCUM_INNER_LOOP_acc_987_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_991_nl = ACCUM_INNER_LOOP_acc_988_nl + ACCUM_INNER_LOOP_acc_987_nl;
  assign ACCUM_INNER_LOOP_acc_991_nl = nl_ACCUM_INNER_LOOP_acc_991_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_992_nl
      + ACCUM_INNER_LOOP_acc_991_nl;
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1 = (ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5349:5345]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5354:5350]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5329:5325]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5334:5330]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5339:5335]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5344:5340]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5359:5355]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5364:5360]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1005_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1005_nl = nl_ACCUM_INNER_LOOP_acc_1005_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5369:5365]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5374:5370]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5379:5375]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5384:5380]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1001_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1001_nl = nl_ACCUM_INNER_LOOP_acc_1001_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1745_nl = (ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[384:380]);
  assign ACCUM_INNER_LOOP_acc_1745_nl = nl_ACCUM_INNER_LOOP_acc_1745_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5324:5320]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1000_nl = ({ACCUM_INNER_LOOP_acc_1745_nl , (ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1000_nl = nl_ACCUM_INNER_LOOP_acc_1000_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1004_nl = ACCUM_INNER_LOOP_acc_1001_nl + ACCUM_INNER_LOOP_acc_1000_nl;
  assign ACCUM_INNER_LOOP_acc_1004_nl = nl_ACCUM_INNER_LOOP_acc_1004_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1005_nl
      + ACCUM_INNER_LOOP_acc_1004_nl;
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1 = (ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5419:5415]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5424:5420]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5399:5395]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5404:5400]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5409:5405]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5414:5410]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5429:5425]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5434:5430]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1018_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1018_nl = nl_ACCUM_INNER_LOOP_acc_1018_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5439:5435]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5444:5440]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5449:5445]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5454:5450]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1014_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1014_nl = nl_ACCUM_INNER_LOOP_acc_1014_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1746_nl = (ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[389:385]);
  assign ACCUM_INNER_LOOP_acc_1746_nl = nl_ACCUM_INNER_LOOP_acc_1746_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5394:5390]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1013_nl = ({ACCUM_INNER_LOOP_acc_1746_nl , (ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1013_nl = nl_ACCUM_INNER_LOOP_acc_1013_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1017_nl = ACCUM_INNER_LOOP_acc_1014_nl + ACCUM_INNER_LOOP_acc_1013_nl;
  assign ACCUM_INNER_LOOP_acc_1017_nl = nl_ACCUM_INNER_LOOP_acc_1017_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1018_nl
      + ACCUM_INNER_LOOP_acc_1017_nl;
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1 = (ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5489:5485]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5494:5490]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5469:5465]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5474:5470]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5479:5475]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5484:5480]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5499:5495]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5504:5500]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1031_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1031_nl = nl_ACCUM_INNER_LOOP_acc_1031_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5509:5505]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5514:5510]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5519:5515]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5524:5520]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1027_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1027_nl = nl_ACCUM_INNER_LOOP_acc_1027_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1747_nl = (ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[394:390]);
  assign ACCUM_INNER_LOOP_acc_1747_nl = nl_ACCUM_INNER_LOOP_acc_1747_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5464:5460]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1026_nl = ({ACCUM_INNER_LOOP_acc_1747_nl , (ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1026_nl = nl_ACCUM_INNER_LOOP_acc_1026_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1030_nl = ACCUM_INNER_LOOP_acc_1027_nl + ACCUM_INNER_LOOP_acc_1026_nl;
  assign ACCUM_INNER_LOOP_acc_1030_nl = nl_ACCUM_INNER_LOOP_acc_1030_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1031_nl
      + ACCUM_INNER_LOOP_acc_1030_nl;
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1 = (ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5559:5555]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5564:5560]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5539:5535]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5544:5540]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5549:5545]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5554:5550]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5569:5565]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5574:5570]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1044_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1044_nl = nl_ACCUM_INNER_LOOP_acc_1044_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5579:5575]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5584:5580]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5589:5585]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5594:5590]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1040_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1040_nl = nl_ACCUM_INNER_LOOP_acc_1040_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1748_nl = (ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[399:395]);
  assign ACCUM_INNER_LOOP_acc_1748_nl = nl_ACCUM_INNER_LOOP_acc_1748_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5534:5530]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1039_nl = ({ACCUM_INNER_LOOP_acc_1748_nl , (ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1039_nl = nl_ACCUM_INNER_LOOP_acc_1039_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1043_nl = ACCUM_INNER_LOOP_acc_1040_nl + ACCUM_INNER_LOOP_acc_1039_nl;
  assign ACCUM_INNER_LOOP_acc_1043_nl = nl_ACCUM_INNER_LOOP_acc_1043_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1044_nl
      + ACCUM_INNER_LOOP_acc_1043_nl;
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1 = (ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5629:5625]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5634:5630]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5609:5605]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5614:5610]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5619:5615]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5624:5620]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5639:5635]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5644:5640]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1057_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1057_nl = nl_ACCUM_INNER_LOOP_acc_1057_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5649:5645]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5654:5650]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5659:5655]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5664:5660]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1053_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1053_nl = nl_ACCUM_INNER_LOOP_acc_1053_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1749_nl = (ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[404:400]);
  assign ACCUM_INNER_LOOP_acc_1749_nl = nl_ACCUM_INNER_LOOP_acc_1749_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5604:5600]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1052_nl = ({ACCUM_INNER_LOOP_acc_1749_nl , (ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1052_nl = nl_ACCUM_INNER_LOOP_acc_1052_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1056_nl = ACCUM_INNER_LOOP_acc_1053_nl + ACCUM_INNER_LOOP_acc_1052_nl;
  assign ACCUM_INNER_LOOP_acc_1056_nl = nl_ACCUM_INNER_LOOP_acc_1056_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1057_nl
      + ACCUM_INNER_LOOP_acc_1056_nl;
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1 = (ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5699:5695]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5704:5700]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5679:5675]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5684:5680]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5689:5685]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5694:5690]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5709:5705]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5714:5710]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1070_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1070_nl = nl_ACCUM_INNER_LOOP_acc_1070_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5719:5715]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5724:5720]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5729:5725]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5734:5730]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1066_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1066_nl = nl_ACCUM_INNER_LOOP_acc_1066_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1750_nl = (ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[409:405]);
  assign ACCUM_INNER_LOOP_acc_1750_nl = nl_ACCUM_INNER_LOOP_acc_1750_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5674:5670]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1065_nl = ({ACCUM_INNER_LOOP_acc_1750_nl , (ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1065_nl = nl_ACCUM_INNER_LOOP_acc_1065_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1069_nl = ACCUM_INNER_LOOP_acc_1066_nl + ACCUM_INNER_LOOP_acc_1065_nl;
  assign ACCUM_INNER_LOOP_acc_1069_nl = nl_ACCUM_INNER_LOOP_acc_1069_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1070_nl
      + ACCUM_INNER_LOOP_acc_1069_nl;
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1 = (ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5769:5765]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5774:5770]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5749:5745]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5754:5750]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5759:5755]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5764:5760]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5779:5775]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5784:5780]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1083_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1083_nl = nl_ACCUM_INNER_LOOP_acc_1083_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5789:5785]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5794:5790]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5799:5795]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5804:5800]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1079_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1079_nl = nl_ACCUM_INNER_LOOP_acc_1079_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1751_nl = (ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[414:410]);
  assign ACCUM_INNER_LOOP_acc_1751_nl = nl_ACCUM_INNER_LOOP_acc_1751_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5744:5740]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1078_nl = ({ACCUM_INNER_LOOP_acc_1751_nl , (ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1078_nl = nl_ACCUM_INNER_LOOP_acc_1078_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1082_nl = ACCUM_INNER_LOOP_acc_1079_nl + ACCUM_INNER_LOOP_acc_1078_nl;
  assign ACCUM_INNER_LOOP_acc_1082_nl = nl_ACCUM_INNER_LOOP_acc_1082_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1083_nl
      + ACCUM_INNER_LOOP_acc_1082_nl;
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1 = (ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5839:5835]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5844:5840]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5819:5815]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5824:5820]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5829:5825]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5834:5830]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5849:5845]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5854:5850]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1096_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1096_nl = nl_ACCUM_INNER_LOOP_acc_1096_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5859:5855]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5864:5860]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5869:5865]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5874:5870]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1092_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1092_nl = nl_ACCUM_INNER_LOOP_acc_1092_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1752_nl = (ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[419:415]);
  assign ACCUM_INNER_LOOP_acc_1752_nl = nl_ACCUM_INNER_LOOP_acc_1752_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5814:5810]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1091_nl = ({ACCUM_INNER_LOOP_acc_1752_nl , (ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1091_nl = nl_ACCUM_INNER_LOOP_acc_1091_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1095_nl = ACCUM_INNER_LOOP_acc_1092_nl + ACCUM_INNER_LOOP_acc_1091_nl;
  assign ACCUM_INNER_LOOP_acc_1095_nl = nl_ACCUM_INNER_LOOP_acc_1095_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1096_nl
      + ACCUM_INNER_LOOP_acc_1095_nl;
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1 = (ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5909:5905]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5914:5910]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5889:5885]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5894:5890]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5899:5895]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5904:5900]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5919:5915]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5924:5920]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1109_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1109_nl = nl_ACCUM_INNER_LOOP_acc_1109_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5929:5925]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[5934:5930]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[5939:5935]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[5944:5940]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1105_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1105_nl = nl_ACCUM_INNER_LOOP_acc_1105_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1753_nl = (ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[424:420]);
  assign ACCUM_INNER_LOOP_acc_1753_nl = nl_ACCUM_INNER_LOOP_acc_1753_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5884:5880]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1104_nl = ({ACCUM_INNER_LOOP_acc_1753_nl , (ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1104_nl = nl_ACCUM_INNER_LOOP_acc_1104_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1108_nl = ACCUM_INNER_LOOP_acc_1105_nl + ACCUM_INNER_LOOP_acc_1104_nl;
  assign ACCUM_INNER_LOOP_acc_1108_nl = nl_ACCUM_INNER_LOOP_acc_1108_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1109_nl
      + ACCUM_INNER_LOOP_acc_1108_nl;
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1 = (ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[5979:5975]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[5984:5980]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[5959:5955]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[5964:5960]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[5969:5965]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[5974:5970]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[5989:5985]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[5994:5990]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1122_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1122_nl = nl_ACCUM_INNER_LOOP_acc_1122_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[5999:5995]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6004:6000]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6009:6005]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6014:6010]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1118_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1118_nl = nl_ACCUM_INNER_LOOP_acc_1118_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1754_nl = (ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[429:425]);
  assign ACCUM_INNER_LOOP_acc_1754_nl = nl_ACCUM_INNER_LOOP_acc_1754_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[5954:5950]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1117_nl = ({ACCUM_INNER_LOOP_acc_1754_nl , (ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1117_nl = nl_ACCUM_INNER_LOOP_acc_1117_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1121_nl = ACCUM_INNER_LOOP_acc_1118_nl + ACCUM_INNER_LOOP_acc_1117_nl;
  assign ACCUM_INNER_LOOP_acc_1121_nl = nl_ACCUM_INNER_LOOP_acc_1121_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1122_nl
      + ACCUM_INNER_LOOP_acc_1121_nl;
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1 = (ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6049:6045]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6054:6050]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6029:6025]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6034:6030]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6039:6035]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6044:6040]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6059:6055]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6064:6060]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1135_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1135_nl = nl_ACCUM_INNER_LOOP_acc_1135_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6069:6065]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6074:6070]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6079:6075]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6084:6080]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1131_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1131_nl = nl_ACCUM_INNER_LOOP_acc_1131_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1755_nl = (ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[434:430]);
  assign ACCUM_INNER_LOOP_acc_1755_nl = nl_ACCUM_INNER_LOOP_acc_1755_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6024:6020]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1130_nl = ({ACCUM_INNER_LOOP_acc_1755_nl , (ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1130_nl = nl_ACCUM_INNER_LOOP_acc_1130_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1134_nl = ACCUM_INNER_LOOP_acc_1131_nl + ACCUM_INNER_LOOP_acc_1130_nl;
  assign ACCUM_INNER_LOOP_acc_1134_nl = nl_ACCUM_INNER_LOOP_acc_1134_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1135_nl
      + ACCUM_INNER_LOOP_acc_1134_nl;
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1 = (ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6119:6115]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6124:6120]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6099:6095]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6104:6100]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6109:6105]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6114:6110]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6129:6125]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6134:6130]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1148_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1148_nl = nl_ACCUM_INNER_LOOP_acc_1148_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6139:6135]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6144:6140]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6149:6145]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6154:6150]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1144_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1144_nl = nl_ACCUM_INNER_LOOP_acc_1144_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1756_nl = (ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[439:435]);
  assign ACCUM_INNER_LOOP_acc_1756_nl = nl_ACCUM_INNER_LOOP_acc_1756_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6094:6090]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1143_nl = ({ACCUM_INNER_LOOP_acc_1756_nl , (ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1143_nl = nl_ACCUM_INNER_LOOP_acc_1143_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1147_nl = ACCUM_INNER_LOOP_acc_1144_nl + ACCUM_INNER_LOOP_acc_1143_nl;
  assign ACCUM_INNER_LOOP_acc_1147_nl = nl_ACCUM_INNER_LOOP_acc_1147_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1148_nl
      + ACCUM_INNER_LOOP_acc_1147_nl;
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1 = (ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6189:6185]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6194:6190]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6169:6165]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6174:6170]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6179:6175]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6184:6180]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6199:6195]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6204:6200]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1161_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1161_nl = nl_ACCUM_INNER_LOOP_acc_1161_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6209:6205]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6214:6210]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6219:6215]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6224:6220]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1157_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1157_nl = nl_ACCUM_INNER_LOOP_acc_1157_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1757_nl = (ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[444:440]);
  assign ACCUM_INNER_LOOP_acc_1757_nl = nl_ACCUM_INNER_LOOP_acc_1757_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6164:6160]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1156_nl = ({ACCUM_INNER_LOOP_acc_1757_nl , (ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1156_nl = nl_ACCUM_INNER_LOOP_acc_1156_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1160_nl = ACCUM_INNER_LOOP_acc_1157_nl + ACCUM_INNER_LOOP_acc_1156_nl;
  assign ACCUM_INNER_LOOP_acc_1160_nl = nl_ACCUM_INNER_LOOP_acc_1160_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1161_nl
      + ACCUM_INNER_LOOP_acc_1160_nl;
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1 = (ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6259:6255]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6264:6260]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6239:6235]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6244:6240]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6249:6245]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6254:6250]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6269:6265]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6274:6270]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1174_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1174_nl = nl_ACCUM_INNER_LOOP_acc_1174_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6279:6275]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6284:6280]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6289:6285]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6294:6290]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1170_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1170_nl = nl_ACCUM_INNER_LOOP_acc_1170_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1758_nl = (ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[449:445]);
  assign ACCUM_INNER_LOOP_acc_1758_nl = nl_ACCUM_INNER_LOOP_acc_1758_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6234:6230]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1169_nl = ({ACCUM_INNER_LOOP_acc_1758_nl , (ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1169_nl = nl_ACCUM_INNER_LOOP_acc_1169_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1173_nl = ACCUM_INNER_LOOP_acc_1170_nl + ACCUM_INNER_LOOP_acc_1169_nl;
  assign ACCUM_INNER_LOOP_acc_1173_nl = nl_ACCUM_INNER_LOOP_acc_1173_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1174_nl
      + ACCUM_INNER_LOOP_acc_1173_nl;
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1 = (ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6329:6325]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6334:6330]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6309:6305]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6314:6310]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6319:6315]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6324:6320]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6339:6335]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6344:6340]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1187_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1187_nl = nl_ACCUM_INNER_LOOP_acc_1187_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6349:6345]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6354:6350]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6359:6355]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6364:6360]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1183_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1183_nl = nl_ACCUM_INNER_LOOP_acc_1183_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1759_nl = (ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[454:450]);
  assign ACCUM_INNER_LOOP_acc_1759_nl = nl_ACCUM_INNER_LOOP_acc_1759_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6304:6300]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1182_nl = ({ACCUM_INNER_LOOP_acc_1759_nl , (ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1182_nl = nl_ACCUM_INNER_LOOP_acc_1182_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1186_nl = ACCUM_INNER_LOOP_acc_1183_nl + ACCUM_INNER_LOOP_acc_1182_nl;
  assign ACCUM_INNER_LOOP_acc_1186_nl = nl_ACCUM_INNER_LOOP_acc_1186_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1187_nl
      + ACCUM_INNER_LOOP_acc_1186_nl;
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1 = (ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6399:6395]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6404:6400]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6379:6375]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6384:6380]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6389:6385]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6394:6390]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6409:6405]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6414:6410]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1200_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1200_nl = nl_ACCUM_INNER_LOOP_acc_1200_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6419:6415]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6424:6420]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6429:6425]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6434:6430]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1196_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1196_nl = nl_ACCUM_INNER_LOOP_acc_1196_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1760_nl = (ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[459:455]);
  assign ACCUM_INNER_LOOP_acc_1760_nl = nl_ACCUM_INNER_LOOP_acc_1760_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6374:6370]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1195_nl = ({ACCUM_INNER_LOOP_acc_1760_nl , (ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1195_nl = nl_ACCUM_INNER_LOOP_acc_1195_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1199_nl = ACCUM_INNER_LOOP_acc_1196_nl + ACCUM_INNER_LOOP_acc_1195_nl;
  assign ACCUM_INNER_LOOP_acc_1199_nl = nl_ACCUM_INNER_LOOP_acc_1199_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1200_nl
      + ACCUM_INNER_LOOP_acc_1199_nl;
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1 = (ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6469:6465]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6474:6470]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6449:6445]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6454:6450]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6459:6455]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6464:6460]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6479:6475]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6484:6480]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1213_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1213_nl = nl_ACCUM_INNER_LOOP_acc_1213_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6489:6485]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6494:6490]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6499:6495]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6504:6500]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1209_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1209_nl = nl_ACCUM_INNER_LOOP_acc_1209_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1761_nl = (ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[464:460]);
  assign ACCUM_INNER_LOOP_acc_1761_nl = nl_ACCUM_INNER_LOOP_acc_1761_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6444:6440]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1208_nl = ({ACCUM_INNER_LOOP_acc_1761_nl , (ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1208_nl = nl_ACCUM_INNER_LOOP_acc_1208_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1212_nl = ACCUM_INNER_LOOP_acc_1209_nl + ACCUM_INNER_LOOP_acc_1208_nl;
  assign ACCUM_INNER_LOOP_acc_1212_nl = nl_ACCUM_INNER_LOOP_acc_1212_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1213_nl
      + ACCUM_INNER_LOOP_acc_1212_nl;
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1 = (ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6539:6535]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6544:6540]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6519:6515]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6524:6520]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6529:6525]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6534:6530]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6549:6545]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6554:6550]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1226_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1226_nl = nl_ACCUM_INNER_LOOP_acc_1226_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6559:6555]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6564:6560]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6569:6565]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6574:6570]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1222_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1222_nl = nl_ACCUM_INNER_LOOP_acc_1222_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1762_nl = (ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[469:465]);
  assign ACCUM_INNER_LOOP_acc_1762_nl = nl_ACCUM_INNER_LOOP_acc_1762_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6514:6510]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1221_nl = ({ACCUM_INNER_LOOP_acc_1762_nl , (ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1221_nl = nl_ACCUM_INNER_LOOP_acc_1221_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1225_nl = ACCUM_INNER_LOOP_acc_1222_nl + ACCUM_INNER_LOOP_acc_1221_nl;
  assign ACCUM_INNER_LOOP_acc_1225_nl = nl_ACCUM_INNER_LOOP_acc_1225_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1226_nl
      + ACCUM_INNER_LOOP_acc_1225_nl;
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1 = (ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6609:6605]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6614:6610]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6589:6585]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6594:6590]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6599:6595]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6604:6600]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6619:6615]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6624:6620]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1239_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1239_nl = nl_ACCUM_INNER_LOOP_acc_1239_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6629:6625]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6634:6630]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6639:6635]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6644:6640]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1235_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1235_nl = nl_ACCUM_INNER_LOOP_acc_1235_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1763_nl = (ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[474:470]);
  assign ACCUM_INNER_LOOP_acc_1763_nl = nl_ACCUM_INNER_LOOP_acc_1763_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6584:6580]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1234_nl = ({ACCUM_INNER_LOOP_acc_1763_nl , (ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1234_nl = nl_ACCUM_INNER_LOOP_acc_1234_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1238_nl = ACCUM_INNER_LOOP_acc_1235_nl + ACCUM_INNER_LOOP_acc_1234_nl;
  assign ACCUM_INNER_LOOP_acc_1238_nl = nl_ACCUM_INNER_LOOP_acc_1238_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1239_nl
      + ACCUM_INNER_LOOP_acc_1238_nl;
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1 = (ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6679:6675]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6684:6680]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6659:6655]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6664:6660]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6669:6665]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6674:6670]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6689:6685]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6694:6690]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1252_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1252_nl = nl_ACCUM_INNER_LOOP_acc_1252_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6699:6695]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6704:6700]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6709:6705]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6714:6710]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1248_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1248_nl = nl_ACCUM_INNER_LOOP_acc_1248_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1764_nl = (ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[479:475]);
  assign ACCUM_INNER_LOOP_acc_1764_nl = nl_ACCUM_INNER_LOOP_acc_1764_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6654:6650]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1247_nl = ({ACCUM_INNER_LOOP_acc_1764_nl , (ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1247_nl = nl_ACCUM_INNER_LOOP_acc_1247_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1251_nl = ACCUM_INNER_LOOP_acc_1248_nl + ACCUM_INNER_LOOP_acc_1247_nl;
  assign ACCUM_INNER_LOOP_acc_1251_nl = nl_ACCUM_INNER_LOOP_acc_1251_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1252_nl
      + ACCUM_INNER_LOOP_acc_1251_nl;
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1 = (ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6749:6745]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6754:6750]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6729:6725]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6734:6730]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6739:6735]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6744:6740]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6759:6755]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6764:6760]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1265_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1265_nl = nl_ACCUM_INNER_LOOP_acc_1265_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6769:6765]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6774:6770]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6779:6775]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6784:6780]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1261_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1261_nl = nl_ACCUM_INNER_LOOP_acc_1261_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1765_nl = (ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[484:480]);
  assign ACCUM_INNER_LOOP_acc_1765_nl = nl_ACCUM_INNER_LOOP_acc_1765_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6724:6720]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1260_nl = ({ACCUM_INNER_LOOP_acc_1765_nl , (ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1260_nl = nl_ACCUM_INNER_LOOP_acc_1260_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1264_nl = ACCUM_INNER_LOOP_acc_1261_nl + ACCUM_INNER_LOOP_acc_1260_nl;
  assign ACCUM_INNER_LOOP_acc_1264_nl = nl_ACCUM_INNER_LOOP_acc_1264_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1265_nl
      + ACCUM_INNER_LOOP_acc_1264_nl;
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1 = (ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6819:6815]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6824:6820]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6799:6795]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6804:6800]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6809:6805]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6814:6810]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6829:6825]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6834:6830]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1278_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1278_nl = nl_ACCUM_INNER_LOOP_acc_1278_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6839:6835]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6844:6840]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6849:6845]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6854:6850]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1274_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1274_nl = nl_ACCUM_INNER_LOOP_acc_1274_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1766_nl = (ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[489:485]);
  assign ACCUM_INNER_LOOP_acc_1766_nl = nl_ACCUM_INNER_LOOP_acc_1766_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6794:6790]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1273_nl = ({ACCUM_INNER_LOOP_acc_1766_nl , (ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1273_nl = nl_ACCUM_INNER_LOOP_acc_1273_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1277_nl = ACCUM_INNER_LOOP_acc_1274_nl + ACCUM_INNER_LOOP_acc_1273_nl;
  assign ACCUM_INNER_LOOP_acc_1277_nl = nl_ACCUM_INNER_LOOP_acc_1277_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1278_nl
      + ACCUM_INNER_LOOP_acc_1277_nl;
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1 = (ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6889:6885]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6894:6890]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6869:6865]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6874:6870]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6879:6875]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6884:6880]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6899:6895]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6904:6900]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1291_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1291_nl = nl_ACCUM_INNER_LOOP_acc_1291_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6909:6905]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6914:6910]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6919:6915]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6924:6920]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1287_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1287_nl = nl_ACCUM_INNER_LOOP_acc_1287_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1767_nl = (ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[494:490]);
  assign ACCUM_INNER_LOOP_acc_1767_nl = nl_ACCUM_INNER_LOOP_acc_1767_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6864:6860]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1286_nl = ({ACCUM_INNER_LOOP_acc_1767_nl , (ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1286_nl = nl_ACCUM_INNER_LOOP_acc_1286_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1290_nl = ACCUM_INNER_LOOP_acc_1287_nl + ACCUM_INNER_LOOP_acc_1286_nl;
  assign ACCUM_INNER_LOOP_acc_1290_nl = nl_ACCUM_INNER_LOOP_acc_1290_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1291_nl
      + ACCUM_INNER_LOOP_acc_1290_nl;
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1 = (ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[6959:6955]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[6964:6960]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[6939:6935]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[6944:6940]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[6949:6945]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[6954:6950]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[6969:6965]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[6974:6970]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1304_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1304_nl = nl_ACCUM_INNER_LOOP_acc_1304_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[6979:6975]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[6984:6980]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[6989:6985]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[6994:6990]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1300_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1300_nl = nl_ACCUM_INNER_LOOP_acc_1300_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1768_nl = (ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[499:495]);
  assign ACCUM_INNER_LOOP_acc_1768_nl = nl_ACCUM_INNER_LOOP_acc_1768_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[6934:6930]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1299_nl = ({ACCUM_INNER_LOOP_acc_1768_nl , (ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1299_nl = nl_ACCUM_INNER_LOOP_acc_1299_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1303_nl = ACCUM_INNER_LOOP_acc_1300_nl + ACCUM_INNER_LOOP_acc_1299_nl;
  assign ACCUM_INNER_LOOP_acc_1303_nl = nl_ACCUM_INNER_LOOP_acc_1303_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1304_nl
      + ACCUM_INNER_LOOP_acc_1303_nl;
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1 = (ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7029:7025]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7034:7030]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7009:7005]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7014:7010]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7019:7015]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7024:7020]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7039:7035]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7044:7040]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1317_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1317_nl = nl_ACCUM_INNER_LOOP_acc_1317_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7049:7045]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7054:7050]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7059:7055]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7064:7060]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1313_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1313_nl = nl_ACCUM_INNER_LOOP_acc_1313_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1769_nl = (ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[504:500]);
  assign ACCUM_INNER_LOOP_acc_1769_nl = nl_ACCUM_INNER_LOOP_acc_1769_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7004:7000]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1312_nl = ({ACCUM_INNER_LOOP_acc_1769_nl , (ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1312_nl = nl_ACCUM_INNER_LOOP_acc_1312_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1316_nl = ACCUM_INNER_LOOP_acc_1313_nl + ACCUM_INNER_LOOP_acc_1312_nl;
  assign ACCUM_INNER_LOOP_acc_1316_nl = nl_ACCUM_INNER_LOOP_acc_1316_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1317_nl
      + ACCUM_INNER_LOOP_acc_1316_nl;
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1 = (ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7099:7095]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7104:7100]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7079:7075]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7084:7080]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7089:7085]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7094:7090]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7109:7105]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7114:7110]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1330_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1330_nl = nl_ACCUM_INNER_LOOP_acc_1330_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7119:7115]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7124:7120]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7129:7125]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7134:7130]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1326_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1326_nl = nl_ACCUM_INNER_LOOP_acc_1326_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1770_nl = (ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[509:505]);
  assign ACCUM_INNER_LOOP_acc_1770_nl = nl_ACCUM_INNER_LOOP_acc_1770_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7074:7070]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1325_nl = ({ACCUM_INNER_LOOP_acc_1770_nl , (ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1325_nl = nl_ACCUM_INNER_LOOP_acc_1325_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1329_nl = ACCUM_INNER_LOOP_acc_1326_nl + ACCUM_INNER_LOOP_acc_1325_nl;
  assign ACCUM_INNER_LOOP_acc_1329_nl = nl_ACCUM_INNER_LOOP_acc_1329_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1330_nl
      + ACCUM_INNER_LOOP_acc_1329_nl;
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1 = (ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7169:7165]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7174:7170]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7149:7145]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7154:7150]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7159:7155]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7164:7160]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7179:7175]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7184:7180]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1343_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1343_nl = nl_ACCUM_INNER_LOOP_acc_1343_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7189:7185]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7194:7190]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7199:7195]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7204:7200]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1339_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1339_nl = nl_ACCUM_INNER_LOOP_acc_1339_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1771_nl = (ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[514:510]);
  assign ACCUM_INNER_LOOP_acc_1771_nl = nl_ACCUM_INNER_LOOP_acc_1771_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7144:7140]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1338_nl = ({ACCUM_INNER_LOOP_acc_1771_nl , (ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1338_nl = nl_ACCUM_INNER_LOOP_acc_1338_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1342_nl = ACCUM_INNER_LOOP_acc_1339_nl + ACCUM_INNER_LOOP_acc_1338_nl;
  assign ACCUM_INNER_LOOP_acc_1342_nl = nl_ACCUM_INNER_LOOP_acc_1342_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1343_nl
      + ACCUM_INNER_LOOP_acc_1342_nl;
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1 = (ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7239:7235]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7244:7240]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7219:7215]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7224:7220]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7229:7225]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7234:7230]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7249:7245]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7254:7250]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1356_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1356_nl = nl_ACCUM_INNER_LOOP_acc_1356_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7259:7255]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7264:7260]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7269:7265]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7274:7270]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1352_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1352_nl = nl_ACCUM_INNER_LOOP_acc_1352_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1772_nl = (ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[519:515]);
  assign ACCUM_INNER_LOOP_acc_1772_nl = nl_ACCUM_INNER_LOOP_acc_1772_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7214:7210]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1351_nl = ({ACCUM_INNER_LOOP_acc_1772_nl , (ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1351_nl = nl_ACCUM_INNER_LOOP_acc_1351_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1355_nl = ACCUM_INNER_LOOP_acc_1352_nl + ACCUM_INNER_LOOP_acc_1351_nl;
  assign ACCUM_INNER_LOOP_acc_1355_nl = nl_ACCUM_INNER_LOOP_acc_1355_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1356_nl
      + ACCUM_INNER_LOOP_acc_1355_nl;
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1 = (ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7309:7305]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7314:7310]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7289:7285]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7294:7290]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7299:7295]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7304:7300]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7319:7315]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7324:7320]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1369_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1369_nl = nl_ACCUM_INNER_LOOP_acc_1369_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7329:7325]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7334:7330]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7339:7335]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7344:7340]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1365_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1365_nl = nl_ACCUM_INNER_LOOP_acc_1365_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1773_nl = (ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[524:520]);
  assign ACCUM_INNER_LOOP_acc_1773_nl = nl_ACCUM_INNER_LOOP_acc_1773_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7284:7280]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1364_nl = ({ACCUM_INNER_LOOP_acc_1773_nl , (ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1364_nl = nl_ACCUM_INNER_LOOP_acc_1364_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1368_nl = ACCUM_INNER_LOOP_acc_1365_nl + ACCUM_INNER_LOOP_acc_1364_nl;
  assign ACCUM_INNER_LOOP_acc_1368_nl = nl_ACCUM_INNER_LOOP_acc_1368_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1369_nl
      + ACCUM_INNER_LOOP_acc_1368_nl;
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1 = (ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7379:7375]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7384:7380]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7359:7355]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7364:7360]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7369:7365]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7374:7370]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7389:7385]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7394:7390]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1382_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1382_nl = nl_ACCUM_INNER_LOOP_acc_1382_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7399:7395]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7404:7400]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7409:7405]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7414:7410]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1378_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1378_nl = nl_ACCUM_INNER_LOOP_acc_1378_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1774_nl = (ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[529:525]);
  assign ACCUM_INNER_LOOP_acc_1774_nl = nl_ACCUM_INNER_LOOP_acc_1774_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7354:7350]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1377_nl = ({ACCUM_INNER_LOOP_acc_1774_nl , (ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1377_nl = nl_ACCUM_INNER_LOOP_acc_1377_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1381_nl = ACCUM_INNER_LOOP_acc_1378_nl + ACCUM_INNER_LOOP_acc_1377_nl;
  assign ACCUM_INNER_LOOP_acc_1381_nl = nl_ACCUM_INNER_LOOP_acc_1381_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1382_nl
      + ACCUM_INNER_LOOP_acc_1381_nl;
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1 = (ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7449:7445]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7454:7450]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7429:7425]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7434:7430]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7439:7435]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7444:7440]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7459:7455]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7464:7460]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1395_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1395_nl = nl_ACCUM_INNER_LOOP_acc_1395_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7469:7465]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7474:7470]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7479:7475]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7484:7480]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1391_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1391_nl = nl_ACCUM_INNER_LOOP_acc_1391_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1775_nl = (ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[534:530]);
  assign ACCUM_INNER_LOOP_acc_1775_nl = nl_ACCUM_INNER_LOOP_acc_1775_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7424:7420]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1390_nl = ({ACCUM_INNER_LOOP_acc_1775_nl , (ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1390_nl = nl_ACCUM_INNER_LOOP_acc_1390_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1394_nl = ACCUM_INNER_LOOP_acc_1391_nl + ACCUM_INNER_LOOP_acc_1390_nl;
  assign ACCUM_INNER_LOOP_acc_1394_nl = nl_ACCUM_INNER_LOOP_acc_1394_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1395_nl
      + ACCUM_INNER_LOOP_acc_1394_nl;
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1 = (ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7519:7515]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7524:7520]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7499:7495]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7504:7500]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7509:7505]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7514:7510]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7529:7525]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7534:7530]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1408_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1408_nl = nl_ACCUM_INNER_LOOP_acc_1408_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7539:7535]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7544:7540]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7549:7545]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7554:7550]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1404_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1404_nl = nl_ACCUM_INNER_LOOP_acc_1404_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1776_nl = (ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[539:535]);
  assign ACCUM_INNER_LOOP_acc_1776_nl = nl_ACCUM_INNER_LOOP_acc_1776_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7494:7490]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1403_nl = ({ACCUM_INNER_LOOP_acc_1776_nl , (ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1403_nl = nl_ACCUM_INNER_LOOP_acc_1403_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1407_nl = ACCUM_INNER_LOOP_acc_1404_nl + ACCUM_INNER_LOOP_acc_1403_nl;
  assign ACCUM_INNER_LOOP_acc_1407_nl = nl_ACCUM_INNER_LOOP_acc_1407_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1408_nl
      + ACCUM_INNER_LOOP_acc_1407_nl;
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1 = (ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7589:7585]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7594:7590]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7569:7565]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7574:7570]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7579:7575]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7584:7580]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7599:7595]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7604:7600]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1421_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1421_nl = nl_ACCUM_INNER_LOOP_acc_1421_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7609:7605]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7614:7610]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7619:7615]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7624:7620]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1417_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1417_nl = nl_ACCUM_INNER_LOOP_acc_1417_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1777_nl = (ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[544:540]);
  assign ACCUM_INNER_LOOP_acc_1777_nl = nl_ACCUM_INNER_LOOP_acc_1777_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7564:7560]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1416_nl = ({ACCUM_INNER_LOOP_acc_1777_nl , (ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1416_nl = nl_ACCUM_INNER_LOOP_acc_1416_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1420_nl = ACCUM_INNER_LOOP_acc_1417_nl + ACCUM_INNER_LOOP_acc_1416_nl;
  assign ACCUM_INNER_LOOP_acc_1420_nl = nl_ACCUM_INNER_LOOP_acc_1420_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1421_nl
      + ACCUM_INNER_LOOP_acc_1420_nl;
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1 = (ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7659:7655]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7664:7660]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7639:7635]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7644:7640]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7649:7645]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7654:7650]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7669:7665]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7674:7670]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1434_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1434_nl = nl_ACCUM_INNER_LOOP_acc_1434_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7679:7675]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7684:7680]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7689:7685]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7694:7690]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1430_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1430_nl = nl_ACCUM_INNER_LOOP_acc_1430_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1778_nl = (ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[549:545]);
  assign ACCUM_INNER_LOOP_acc_1778_nl = nl_ACCUM_INNER_LOOP_acc_1778_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7634:7630]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1429_nl = ({ACCUM_INNER_LOOP_acc_1778_nl , (ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1429_nl = nl_ACCUM_INNER_LOOP_acc_1429_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1433_nl = ACCUM_INNER_LOOP_acc_1430_nl + ACCUM_INNER_LOOP_acc_1429_nl;
  assign ACCUM_INNER_LOOP_acc_1433_nl = nl_ACCUM_INNER_LOOP_acc_1433_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1434_nl
      + ACCUM_INNER_LOOP_acc_1433_nl;
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1 = (ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7729:7725]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7734:7730]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7709:7705]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7714:7710]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7719:7715]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7724:7720]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7739:7735]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7744:7740]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1447_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1447_nl = nl_ACCUM_INNER_LOOP_acc_1447_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7749:7745]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7754:7750]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7759:7755]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7764:7760]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1443_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1443_nl = nl_ACCUM_INNER_LOOP_acc_1443_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1779_nl = (ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[554:550]);
  assign ACCUM_INNER_LOOP_acc_1779_nl = nl_ACCUM_INNER_LOOP_acc_1779_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7704:7700]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1442_nl = ({ACCUM_INNER_LOOP_acc_1779_nl , (ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1442_nl = nl_ACCUM_INNER_LOOP_acc_1442_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1446_nl = ACCUM_INNER_LOOP_acc_1443_nl + ACCUM_INNER_LOOP_acc_1442_nl;
  assign ACCUM_INNER_LOOP_acc_1446_nl = nl_ACCUM_INNER_LOOP_acc_1446_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1447_nl
      + ACCUM_INNER_LOOP_acc_1446_nl;
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1 = (ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7799:7795]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7804:7800]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7779:7775]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7784:7780]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7789:7785]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7794:7790]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7809:7805]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7814:7810]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1460_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1460_nl = nl_ACCUM_INNER_LOOP_acc_1460_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7819:7815]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7824:7820]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7829:7825]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7834:7830]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1456_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1456_nl = nl_ACCUM_INNER_LOOP_acc_1456_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1780_nl = (ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[559:555]);
  assign ACCUM_INNER_LOOP_acc_1780_nl = nl_ACCUM_INNER_LOOP_acc_1780_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7774:7770]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1455_nl = ({ACCUM_INNER_LOOP_acc_1780_nl , (ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1455_nl = nl_ACCUM_INNER_LOOP_acc_1455_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1459_nl = ACCUM_INNER_LOOP_acc_1456_nl + ACCUM_INNER_LOOP_acc_1455_nl;
  assign ACCUM_INNER_LOOP_acc_1459_nl = nl_ACCUM_INNER_LOOP_acc_1459_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1460_nl
      + ACCUM_INNER_LOOP_acc_1459_nl;
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1 = (ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7869:7865]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7874:7870]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7849:7845]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7854:7850]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7859:7855]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7864:7860]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7879:7875]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7884:7880]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1473_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1473_nl = nl_ACCUM_INNER_LOOP_acc_1473_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7889:7885]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7894:7890]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7899:7895]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7904:7900]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1469_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1469_nl = nl_ACCUM_INNER_LOOP_acc_1469_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1781_nl = (ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[564:560]);
  assign ACCUM_INNER_LOOP_acc_1781_nl = nl_ACCUM_INNER_LOOP_acc_1781_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7844:7840]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1468_nl = ({ACCUM_INNER_LOOP_acc_1781_nl , (ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1468_nl = nl_ACCUM_INNER_LOOP_acc_1468_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1472_nl = ACCUM_INNER_LOOP_acc_1469_nl + ACCUM_INNER_LOOP_acc_1468_nl;
  assign ACCUM_INNER_LOOP_acc_1472_nl = nl_ACCUM_INNER_LOOP_acc_1472_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1473_nl
      + ACCUM_INNER_LOOP_acc_1472_nl;
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1 = (ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[7939:7935]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[7944:7940]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7919:7915]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7924:7920]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7929:7925]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[7934:7930]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[7949:7945]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[7954:7950]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1486_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1486_nl = nl_ACCUM_INNER_LOOP_acc_1486_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[7959:7955]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[7964:7960]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[7969:7965]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[7974:7970]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1482_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1482_nl = nl_ACCUM_INNER_LOOP_acc_1482_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1782_nl = (ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[569:565]);
  assign ACCUM_INNER_LOOP_acc_1782_nl = nl_ACCUM_INNER_LOOP_acc_1782_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7914:7910]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1481_nl = ({ACCUM_INNER_LOOP_acc_1782_nl , (ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1481_nl = nl_ACCUM_INNER_LOOP_acc_1481_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1485_nl = ACCUM_INNER_LOOP_acc_1482_nl + ACCUM_INNER_LOOP_acc_1481_nl;
  assign ACCUM_INNER_LOOP_acc_1485_nl = nl_ACCUM_INNER_LOOP_acc_1485_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1486_nl
      + ACCUM_INNER_LOOP_acc_1485_nl;
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1 = (ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8009:8005]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8014:8010]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[7989:7985]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[7994:7990]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[7999:7995]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8004:8000]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8019:8015]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8024:8020]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1499_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1499_nl = nl_ACCUM_INNER_LOOP_acc_1499_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8029:8025]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8034:8030]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8039:8035]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8044:8040]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1495_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1495_nl = nl_ACCUM_INNER_LOOP_acc_1495_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1783_nl = (ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[574:570]);
  assign ACCUM_INNER_LOOP_acc_1783_nl = nl_ACCUM_INNER_LOOP_acc_1783_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[7984:7980]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1494_nl = ({ACCUM_INNER_LOOP_acc_1783_nl , (ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1494_nl = nl_ACCUM_INNER_LOOP_acc_1494_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1498_nl = ACCUM_INNER_LOOP_acc_1495_nl + ACCUM_INNER_LOOP_acc_1494_nl;
  assign ACCUM_INNER_LOOP_acc_1498_nl = nl_ACCUM_INNER_LOOP_acc_1498_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1499_nl
      + ACCUM_INNER_LOOP_acc_1498_nl;
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1 = (ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8079:8075]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8084:8080]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8059:8055]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8064:8060]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8069:8065]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8074:8070]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8089:8085]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8094:8090]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1512_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1512_nl = nl_ACCUM_INNER_LOOP_acc_1512_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8099:8095]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8104:8100]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8109:8105]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8114:8110]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1508_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1508_nl = nl_ACCUM_INNER_LOOP_acc_1508_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1784_nl = (ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[579:575]);
  assign ACCUM_INNER_LOOP_acc_1784_nl = nl_ACCUM_INNER_LOOP_acc_1784_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8054:8050]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1507_nl = ({ACCUM_INNER_LOOP_acc_1784_nl , (ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1507_nl = nl_ACCUM_INNER_LOOP_acc_1507_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1511_nl = ACCUM_INNER_LOOP_acc_1508_nl + ACCUM_INNER_LOOP_acc_1507_nl;
  assign ACCUM_INNER_LOOP_acc_1511_nl = nl_ACCUM_INNER_LOOP_acc_1511_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1512_nl
      + ACCUM_INNER_LOOP_acc_1511_nl;
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1 = (ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8149:8145]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8154:8150]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8129:8125]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8134:8130]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8139:8135]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8144:8140]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8159:8155]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8164:8160]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1525_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1525_nl = nl_ACCUM_INNER_LOOP_acc_1525_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8169:8165]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8174:8170]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8179:8175]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8184:8180]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1521_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1521_nl = nl_ACCUM_INNER_LOOP_acc_1521_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1785_nl = (ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[584:580]);
  assign ACCUM_INNER_LOOP_acc_1785_nl = nl_ACCUM_INNER_LOOP_acc_1785_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8124:8120]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1520_nl = ({ACCUM_INNER_LOOP_acc_1785_nl , (ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1520_nl = nl_ACCUM_INNER_LOOP_acc_1520_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1524_nl = ACCUM_INNER_LOOP_acc_1521_nl + ACCUM_INNER_LOOP_acc_1520_nl;
  assign ACCUM_INNER_LOOP_acc_1524_nl = nl_ACCUM_INNER_LOOP_acc_1524_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1525_nl
      + ACCUM_INNER_LOOP_acc_1524_nl;
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1 = (ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8219:8215]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8224:8220]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8199:8195]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8204:8200]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8209:8205]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8214:8210]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8229:8225]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8234:8230]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1538_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1538_nl = nl_ACCUM_INNER_LOOP_acc_1538_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8239:8235]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8244:8240]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8249:8245]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8254:8250]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1534_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1534_nl = nl_ACCUM_INNER_LOOP_acc_1534_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1786_nl = (ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[589:585]);
  assign ACCUM_INNER_LOOP_acc_1786_nl = nl_ACCUM_INNER_LOOP_acc_1786_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8194:8190]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1533_nl = ({ACCUM_INNER_LOOP_acc_1786_nl , (ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1533_nl = nl_ACCUM_INNER_LOOP_acc_1533_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1537_nl = ACCUM_INNER_LOOP_acc_1534_nl + ACCUM_INNER_LOOP_acc_1533_nl;
  assign ACCUM_INNER_LOOP_acc_1537_nl = nl_ACCUM_INNER_LOOP_acc_1537_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1538_nl
      + ACCUM_INNER_LOOP_acc_1537_nl;
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1 = (ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8289:8285]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8294:8290]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8269:8265]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8274:8270]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8279:8275]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8284:8280]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8299:8295]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8304:8300]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1551_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1551_nl = nl_ACCUM_INNER_LOOP_acc_1551_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8309:8305]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8314:8310]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8319:8315]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8324:8320]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1547_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1547_nl = nl_ACCUM_INNER_LOOP_acc_1547_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1787_nl = (ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[594:590]);
  assign ACCUM_INNER_LOOP_acc_1787_nl = nl_ACCUM_INNER_LOOP_acc_1787_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8264:8260]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1546_nl = ({ACCUM_INNER_LOOP_acc_1787_nl , (ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1546_nl = nl_ACCUM_INNER_LOOP_acc_1546_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1550_nl = ACCUM_INNER_LOOP_acc_1547_nl + ACCUM_INNER_LOOP_acc_1546_nl;
  assign ACCUM_INNER_LOOP_acc_1550_nl = nl_ACCUM_INNER_LOOP_acc_1550_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1551_nl
      + ACCUM_INNER_LOOP_acc_1550_nl;
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1 = (ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8359:8355]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8364:8360]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8339:8335]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8344:8340]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8349:8345]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8354:8350]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8369:8365]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8374:8370]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1564_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1564_nl = nl_ACCUM_INNER_LOOP_acc_1564_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8379:8375]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8384:8380]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8389:8385]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8394:8390]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1560_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1560_nl = nl_ACCUM_INNER_LOOP_acc_1560_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1788_nl = (ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[599:595]);
  assign ACCUM_INNER_LOOP_acc_1788_nl = nl_ACCUM_INNER_LOOP_acc_1788_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8334:8330]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1559_nl = ({ACCUM_INNER_LOOP_acc_1788_nl , (ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1559_nl = nl_ACCUM_INNER_LOOP_acc_1559_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1563_nl = ACCUM_INNER_LOOP_acc_1560_nl + ACCUM_INNER_LOOP_acc_1559_nl;
  assign ACCUM_INNER_LOOP_acc_1563_nl = nl_ACCUM_INNER_LOOP_acc_1563_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1564_nl
      + ACCUM_INNER_LOOP_acc_1563_nl;
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1 = (ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8429:8425]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8434:8430]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8409:8405]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8414:8410]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8419:8415]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8424:8420]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8439:8435]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8444:8440]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1577_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1577_nl = nl_ACCUM_INNER_LOOP_acc_1577_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8449:8445]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8454:8450]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8459:8455]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8464:8460]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1573_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1573_nl = nl_ACCUM_INNER_LOOP_acc_1573_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1789_nl = (ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[604:600]);
  assign ACCUM_INNER_LOOP_acc_1789_nl = nl_ACCUM_INNER_LOOP_acc_1789_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8404:8400]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1572_nl = ({ACCUM_INNER_LOOP_acc_1789_nl , (ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1572_nl = nl_ACCUM_INNER_LOOP_acc_1572_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1576_nl = ACCUM_INNER_LOOP_acc_1573_nl + ACCUM_INNER_LOOP_acc_1572_nl;
  assign ACCUM_INNER_LOOP_acc_1576_nl = nl_ACCUM_INNER_LOOP_acc_1576_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1577_nl
      + ACCUM_INNER_LOOP_acc_1576_nl;
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1 = (ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8499:8495]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8504:8500]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8479:8475]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8484:8480]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8489:8485]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8494:8490]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8509:8505]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8514:8510]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1590_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1590_nl = nl_ACCUM_INNER_LOOP_acc_1590_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8519:8515]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8524:8520]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8529:8525]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8534:8530]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1586_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1586_nl = nl_ACCUM_INNER_LOOP_acc_1586_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1790_nl = (ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[609:605]);
  assign ACCUM_INNER_LOOP_acc_1790_nl = nl_ACCUM_INNER_LOOP_acc_1790_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8474:8470]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1585_nl = ({ACCUM_INNER_LOOP_acc_1790_nl , (ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1585_nl = nl_ACCUM_INNER_LOOP_acc_1585_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1589_nl = ACCUM_INNER_LOOP_acc_1586_nl + ACCUM_INNER_LOOP_acc_1585_nl;
  assign ACCUM_INNER_LOOP_acc_1589_nl = nl_ACCUM_INNER_LOOP_acc_1589_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1590_nl
      + ACCUM_INNER_LOOP_acc_1589_nl;
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1 = (ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8569:8565]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8574:8570]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8549:8545]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8554:8550]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8559:8555]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8564:8560]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8579:8575]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8584:8580]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1603_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1603_nl = nl_ACCUM_INNER_LOOP_acc_1603_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8589:8585]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8594:8590]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8599:8595]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8604:8600]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1599_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1599_nl = nl_ACCUM_INNER_LOOP_acc_1599_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1791_nl = (ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[614:610]);
  assign ACCUM_INNER_LOOP_acc_1791_nl = nl_ACCUM_INNER_LOOP_acc_1791_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8544:8540]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1598_nl = ({ACCUM_INNER_LOOP_acc_1791_nl , (ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1598_nl = nl_ACCUM_INNER_LOOP_acc_1598_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1602_nl = ACCUM_INNER_LOOP_acc_1599_nl + ACCUM_INNER_LOOP_acc_1598_nl;
  assign ACCUM_INNER_LOOP_acc_1602_nl = nl_ACCUM_INNER_LOOP_acc_1602_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1603_nl
      + ACCUM_INNER_LOOP_acc_1602_nl;
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1 = (ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8639:8635]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8644:8640]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8619:8615]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8624:8620]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8629:8625]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8634:8630]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8649:8645]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8654:8650]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1616_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1616_nl = nl_ACCUM_INNER_LOOP_acc_1616_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8659:8655]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8664:8660]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8669:8665]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8674:8670]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1612_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1612_nl = nl_ACCUM_INNER_LOOP_acc_1612_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1792_nl = (ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[619:615]);
  assign ACCUM_INNER_LOOP_acc_1792_nl = nl_ACCUM_INNER_LOOP_acc_1792_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8614:8610]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1611_nl = ({ACCUM_INNER_LOOP_acc_1792_nl , (ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1611_nl = nl_ACCUM_INNER_LOOP_acc_1611_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1615_nl = ACCUM_INNER_LOOP_acc_1612_nl + ACCUM_INNER_LOOP_acc_1611_nl;
  assign ACCUM_INNER_LOOP_acc_1615_nl = nl_ACCUM_INNER_LOOP_acc_1615_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1616_nl
      + ACCUM_INNER_LOOP_acc_1615_nl;
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1 = (ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8709:8705]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8714:8710]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8689:8685]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8694:8690]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8699:8695]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8704:8700]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8719:8715]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8724:8720]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1629_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1629_nl = nl_ACCUM_INNER_LOOP_acc_1629_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8729:8725]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8734:8730]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8739:8735]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8744:8740]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1625_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1625_nl = nl_ACCUM_INNER_LOOP_acc_1625_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1793_nl = (ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[624:620]);
  assign ACCUM_INNER_LOOP_acc_1793_nl = nl_ACCUM_INNER_LOOP_acc_1793_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8684:8680]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1624_nl = ({ACCUM_INNER_LOOP_acc_1793_nl , (ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1624_nl = nl_ACCUM_INNER_LOOP_acc_1624_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1628_nl = ACCUM_INNER_LOOP_acc_1625_nl + ACCUM_INNER_LOOP_acc_1624_nl;
  assign ACCUM_INNER_LOOP_acc_1628_nl = nl_ACCUM_INNER_LOOP_acc_1628_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1629_nl
      + ACCUM_INNER_LOOP_acc_1628_nl;
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1 = (ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8779:8775]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8784:8780]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8759:8755]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8764:8760]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8769:8765]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8774:8770]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8789:8785]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8794:8790]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1642_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1642_nl = nl_ACCUM_INNER_LOOP_acc_1642_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8799:8795]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8804:8800]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8809:8805]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8814:8810]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1638_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1638_nl = nl_ACCUM_INNER_LOOP_acc_1638_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1794_nl = (ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[629:625]);
  assign ACCUM_INNER_LOOP_acc_1794_nl = nl_ACCUM_INNER_LOOP_acc_1794_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8754:8750]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1637_nl = ({ACCUM_INNER_LOOP_acc_1794_nl , (ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1637_nl = nl_ACCUM_INNER_LOOP_acc_1637_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1641_nl = ACCUM_INNER_LOOP_acc_1638_nl + ACCUM_INNER_LOOP_acc_1637_nl;
  assign ACCUM_INNER_LOOP_acc_1641_nl = nl_ACCUM_INNER_LOOP_acc_1641_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1642_nl
      + ACCUM_INNER_LOOP_acc_1641_nl;
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1 = (ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8849:8845]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8854:8850]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8829:8825]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8834:8830]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8839:8835]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8844:8840]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8859:8855]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8864:8860]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1655_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1655_nl = nl_ACCUM_INNER_LOOP_acc_1655_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8869:8865]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8874:8870]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8879:8875]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8884:8880]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1651_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1651_nl = nl_ACCUM_INNER_LOOP_acc_1651_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1795_nl = (ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[634:630]);
  assign ACCUM_INNER_LOOP_acc_1795_nl = nl_ACCUM_INNER_LOOP_acc_1795_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8824:8820]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1650_nl = ({ACCUM_INNER_LOOP_acc_1795_nl , (ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1650_nl = nl_ACCUM_INNER_LOOP_acc_1650_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1654_nl = ACCUM_INNER_LOOP_acc_1651_nl + ACCUM_INNER_LOOP_acc_1650_nl;
  assign ACCUM_INNER_LOOP_acc_1654_nl = nl_ACCUM_INNER_LOOP_acc_1654_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1655_nl
      + ACCUM_INNER_LOOP_acc_1654_nl;
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 = (ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[14:10]!=5'b00000);
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[95:80]))
      * $signed((w2_rsci_idat[8919:8915]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[111:96]))
      * $signed((w2_rsci_idat[8924:8920]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[31:16]))
      * $signed((w2_rsci_idat[8899:8895]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[47:32]))
      * $signed((w2_rsci_idat[8904:8900]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[63:48]))
      * $signed((w2_rsci_idat[8909:8905]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[79:64]))
      * $signed((w2_rsci_idat[8914:8910]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[127:112]))
      * $signed((w2_rsci_idat[8929:8925]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[143:128]))
      * $signed((w2_rsci_idat[8934:8930]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1668_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_6_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_7_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_2_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_3_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_4_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_5_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_8_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_9_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1668_nl = nl_ACCUM_INNER_LOOP_acc_1668_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[159:144]))
      * $signed((w2_rsci_idat[8939:8935]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[175:160]))
      * $signed((w2_rsci_idat[8944:8940]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[191:176]))
      * $signed((w2_rsci_idat[8949:8945]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[207:192]))
      * $signed((w2_rsci_idat[8954:8950]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1664_nl = (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_10_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_11_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_12_ACCUM_INNER_LOOP_mul_nl))
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_13_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1664_nl = nl_ACCUM_INNER_LOOP_acc_1664_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1796_nl = (ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[15:6])
      + conv_s2s_5_10(b2_rsci_idat[639:635]);
  assign ACCUM_INNER_LOOP_acc_1796_nl = nl_ACCUM_INNER_LOOP_acc_1796_nl[9:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[15:0]))
      * $signed((w2_rsci_idat[8894:8890]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign nl_ACCUM_INNER_LOOP_acc_1663_nl = ({ACCUM_INNER_LOOP_acc_1796_nl , (ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1[5:0])})
      + (readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_1_ACCUM_INNER_LOOP_mul_nl));
  assign ACCUM_INNER_LOOP_acc_1663_nl = nl_ACCUM_INNER_LOOP_acc_1663_nl[15:0];
  assign nl_ACCUM_INNER_LOOP_acc_1667_nl = ACCUM_INNER_LOOP_acc_1664_nl + ACCUM_INNER_LOOP_acc_1663_nl;
  assign ACCUM_INNER_LOOP_acc_1667_nl = nl_ACCUM_INNER_LOOP_acc_1667_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = ACCUM_INNER_LOOP_acc_1668_nl
      + ACCUM_INNER_LOOP_acc_1667_nl;
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1 = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_319_9 , layer4_out_conc_319_8_1 , layer4_out_conc_319_0}))
      * $signed((w5_rsci_idat[1289:1285]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1
      = readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_319_9 , layer4_out_conc_319_8_1 , layer4_out_conc_319_0}))
      * $signed((w5_rsci_idat[9:5]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1
      = readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_319_9 , layer4_out_conc_319_8_1 , layer4_out_conc_319_0}))
      * $signed((w5_rsci_idat[649:645]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1
      = readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_16_17(layer2_out_0_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1
      = readslicef_17_1_16(nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8959:8955]));
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8889:8885]));
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8819:8815]));
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8749:8745]));
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8679:8675]));
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8609:8605]));
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8539:8535]));
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8469:8465]));
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8399:8395]));
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8329:8325]));
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8259:8255]));
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8189:8185]));
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8119:8115]));
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[8049:8045]));
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7979:7975]));
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7909:7905]));
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7839:7835]));
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7769:7765]));
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7699:7695]));
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7629:7625]));
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7559:7555]));
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7489:7485]));
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7419:7415]));
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7349:7345]));
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7279:7275]));
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7209:7205]));
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7139:7135]));
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[7069:7065]));
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6999:6995]));
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6929:6925]));
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6859:6855]));
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6789:6785]));
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6719:6715]));
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6649:6645]));
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6579:6575]));
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6509:6505]));
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6439:6435]));
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6369:6365]));
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6299:6295]));
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6229:6225]));
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6159:6155]));
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6089:6085]));
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[6019:6015]));
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5949:5945]));
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5879:5875]));
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5809:5805]));
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5739:5735]));
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5669:5665]));
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5599:5595]));
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5529:5525]));
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5459:5455]));
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5389:5385]));
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5319:5315]));
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5249:5245]));
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5179:5175]));
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5109:5105]));
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[5039:5035]));
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4969:4965]));
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4899:4895]));
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4829:4825]));
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4759:4755]));
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4689:4685]));
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4619:4615]));
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4549:4545]));
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4479:4475]));
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4409:4405]));
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4339:4335]));
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4269:4265]));
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4199:4195]));
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4129:4125]));
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[4059:4055]));
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3989:3985]));
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3919:3915]));
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3849:3845]));
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3779:3775]));
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3709:3705]));
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3639:3635]));
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3569:3565]));
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3499:3495]));
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3429:3425]));
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3359:3355]));
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3289:3285]));
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3219:3215]));
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3149:3145]));
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3079:3075]));
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[3009:3005]));
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2939:2935]));
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2869:2865]));
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2799:2795]));
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2729:2725]));
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2659:2655]));
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2589:2585]));
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2519:2515]));
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2449:2445]));
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2379:2375]));
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2309:2305]));
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2239:2235]));
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2169:2165]));
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2099:2095]));
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[2029:2025]));
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1959:1955]));
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1889:1885]));
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1819:1815]));
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1749:1745]));
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1679:1675]));
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1609:1605]));
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1539:1535]));
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1469:1465]));
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1399:1395]));
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1329:1325]));
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1259:1255]));
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1189:1185]));
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1119:1115]));
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[1049:1045]));
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[979:975]));
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[909:905]));
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[839:835]));
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[769:765]));
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[699:695]));
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1
      = readslicef_20_16_4(ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[629:625]));
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[559:555]));
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[489:485]));
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[419:415]));
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[349:345]));
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[279:275]));
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[209:205]));
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[139:135]));
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = $signed((input_1_rsci_idat[223:208]))
      * $signed((w2_rsci_idat[69:65]));
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl = nl_ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl[19:0];
  assign ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_itm_19_4_1 =
      readslicef_20_16_4(ACCUM_OUTER_LOOP_1_ACCUM_INNER_LOOP_14_ACCUM_INNER_LOOP_mul_nl);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_9 = ((ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_127_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_0 = ((ACCUM_OUTER_LOOP_127_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_127_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_127_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_9 = ((ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_128_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_0 = ((ACCUM_OUTER_LOOP_128_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_128_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_9 = ((ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_125_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_0 = ((ACCUM_OUTER_LOOP_125_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_125_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_125_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_9 = ((ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_126_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_0 = ((ACCUM_OUTER_LOOP_126_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_126_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_126_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_9 = ((ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_123_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_0 = ((ACCUM_OUTER_LOOP_123_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_123_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_123_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_9 = ((ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_124_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_0 = ((ACCUM_OUTER_LOOP_124_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_124_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_124_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_9 = ((ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_121_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_0 = ((ACCUM_OUTER_LOOP_121_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_121_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_121_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_9 = ((ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_122_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_0 = ((ACCUM_OUTER_LOOP_122_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_122_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_122_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_9 = ((ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_119_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_0 = ((ACCUM_OUTER_LOOP_119_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_119_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_119_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_9 = ((ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_120_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_0 = ((ACCUM_OUTER_LOOP_120_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_120_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_120_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_9 = ((ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_117_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_0 = ((ACCUM_OUTER_LOOP_117_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_117_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_117_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_9 = ((ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_118_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_0 = ((ACCUM_OUTER_LOOP_118_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_118_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_118_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_9 = ((ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_115_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_0 = ((ACCUM_OUTER_LOOP_115_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_115_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_115_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_9 = ((ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_116_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_0 = ((ACCUM_OUTER_LOOP_116_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_116_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_116_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_9 = ((ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_113_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_0 = ((ACCUM_OUTER_LOOP_113_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_113_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_113_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_9 = ((ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_114_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_0 = ((ACCUM_OUTER_LOOP_114_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_114_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_114_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_9 = ((ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_111_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_0 = ((ACCUM_OUTER_LOOP_111_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_111_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_111_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_9 = ((ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_112_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_0 = ((ACCUM_OUTER_LOOP_112_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_112_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_112_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_9 = ((ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_109_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_0 = ((ACCUM_OUTER_LOOP_109_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_109_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_109_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_9 = ((ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_110_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_0 = ((ACCUM_OUTER_LOOP_110_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_110_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_110_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_9 = ((ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_107_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_0 = ((ACCUM_OUTER_LOOP_107_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_107_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_107_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_9 = ((ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_108_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_0 = ((ACCUM_OUTER_LOOP_108_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_108_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_108_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_9 = ((ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_105_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_0 = ((ACCUM_OUTER_LOOP_105_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_105_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_105_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_9 = ((ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_106_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_0 = ((ACCUM_OUTER_LOOP_106_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_106_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_106_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_9 = ((ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_103_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_0 = ((ACCUM_OUTER_LOOP_103_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_103_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_103_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_9 = ((ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_104_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_0 = ((ACCUM_OUTER_LOOP_104_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_104_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_104_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_9 = ((ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_101_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_0 = ((ACCUM_OUTER_LOOP_101_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_101_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_101_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_9 = ((ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_102_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_0 = ((ACCUM_OUTER_LOOP_102_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_102_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_102_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_9 = ((ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_99_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_0 = ((ACCUM_OUTER_LOOP_99_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_99_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_99_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_9 = ((ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_100_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_0 = ((ACCUM_OUTER_LOOP_100_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_100_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_100_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_9 = ((ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_97_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_0 = ((ACCUM_OUTER_LOOP_97_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_97_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_97_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_9 = ((ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_98_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_0 = ((ACCUM_OUTER_LOOP_98_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_98_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_98_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_9 = ((ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_95_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_0 = ((ACCUM_OUTER_LOOP_95_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_95_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_95_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_9 = ((ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_96_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_0 = ((ACCUM_OUTER_LOOP_96_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_96_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_96_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_9 = ((ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_93_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_0 = ((ACCUM_OUTER_LOOP_93_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_93_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_93_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_9 = ((ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_94_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_0 = ((ACCUM_OUTER_LOOP_94_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_94_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_94_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_9 = ((ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_91_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_0 = ((ACCUM_OUTER_LOOP_91_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_91_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_91_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_9 = ((ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_92_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_0 = ((ACCUM_OUTER_LOOP_92_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_92_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_92_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_9 = ((ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_89_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_0 = ((ACCUM_OUTER_LOOP_89_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_89_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_89_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_9 = ((ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_90_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_0 = ((ACCUM_OUTER_LOOP_90_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_90_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_90_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_9 = ((ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_87_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_0 = ((ACCUM_OUTER_LOOP_87_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_87_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_87_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_9 = ((ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_88_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_0 = ((ACCUM_OUTER_LOOP_88_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_88_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_88_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_9 = ((ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_85_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_0 = ((ACCUM_OUTER_LOOP_85_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_85_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_85_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_9 = ((ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_86_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_0 = ((ACCUM_OUTER_LOOP_86_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_86_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_86_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_9 = ((ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_83_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_0 = ((ACCUM_OUTER_LOOP_83_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_83_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_83_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_9 = ((ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_84_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_0 = ((ACCUM_OUTER_LOOP_84_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_84_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_84_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_9 = ((ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_81_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_0 = ((ACCUM_OUTER_LOOP_81_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_81_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_81_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_9 = ((ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_82_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_0 = ((ACCUM_OUTER_LOOP_82_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_82_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_82_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_9 = ((ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_79_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_0 = ((ACCUM_OUTER_LOOP_79_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_79_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_79_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_9 = ((ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_80_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_0 = ((ACCUM_OUTER_LOOP_80_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_80_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_80_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_9 = ((ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_77_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_0 = ((ACCUM_OUTER_LOOP_77_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_77_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_77_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_9 = ((ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_78_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_0 = ((ACCUM_OUTER_LOOP_78_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_78_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_78_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_9 = ((ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_75_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_0 = ((ACCUM_OUTER_LOOP_75_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_75_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_75_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_9 = ((ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_76_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_0 = ((ACCUM_OUTER_LOOP_76_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_76_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_76_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_9 = ((ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_73_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_0 = ((ACCUM_OUTER_LOOP_73_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_73_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_73_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_9 = ((ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_74_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_0 = ((ACCUM_OUTER_LOOP_74_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_74_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_74_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_9 = ((ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_71_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_0 = ((ACCUM_OUTER_LOOP_71_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_71_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_71_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_9 = ((ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_72_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_0 = ((ACCUM_OUTER_LOOP_72_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_72_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_72_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_9 = ((ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_69_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_0 = ((ACCUM_OUTER_LOOP_69_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_69_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_69_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_9 = ((ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_70_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_0 = ((ACCUM_OUTER_LOOP_70_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_70_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_70_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_9 = ((ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_67_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_0 = ((ACCUM_OUTER_LOOP_67_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_67_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_67_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_9 = ((ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_68_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_0 = ((ACCUM_OUTER_LOOP_68_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_68_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_68_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_9 = ((ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_65_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_0 = ((ACCUM_OUTER_LOOP_65_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_65_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_65_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_9 = ((ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_8_1 = MUX_v_8_2_2(8'b00000000,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_66_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_0 = ((ACCUM_OUTER_LOOP_66_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_66_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_66_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_193_9 = ((ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1);
  assign layer4_out_conc_193_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_193_0 = ((ACCUM_OUTER_LOOP_63_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_63_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_195_9 = ((ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1);
  assign layer4_out_conc_195_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_195_0 = ((ACCUM_OUTER_LOOP_64_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_64_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_64_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_197_9 = ((ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1);
  assign layer4_out_conc_197_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_197_0 = ((ACCUM_OUTER_LOOP_61_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_61_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_199_9 = ((ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1);
  assign layer4_out_conc_199_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_199_0 = ((ACCUM_OUTER_LOOP_62_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_62_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_201_9 = ((ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1);
  assign layer4_out_conc_201_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_201_0 = ((ACCUM_OUTER_LOOP_59_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_59_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_203_9 = ((ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1);
  assign layer4_out_conc_203_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_203_0 = ((ACCUM_OUTER_LOOP_60_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_60_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_205_9 = ((ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1);
  assign layer4_out_conc_205_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_205_0 = ((ACCUM_OUTER_LOOP_57_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_57_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_207_9 = ((ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1);
  assign layer4_out_conc_207_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_207_0 = ((ACCUM_OUTER_LOOP_58_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_58_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_209_9 = ((ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1);
  assign layer4_out_conc_209_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_209_0 = ((ACCUM_OUTER_LOOP_55_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_55_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_211_9 = ((ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1);
  assign layer4_out_conc_211_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_211_0 = ((ACCUM_OUTER_LOOP_56_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_56_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_213_9 = ((ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1);
  assign layer4_out_conc_213_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_213_0 = ((ACCUM_OUTER_LOOP_53_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_53_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_215_9 = ((ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1);
  assign layer4_out_conc_215_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_215_0 = ((ACCUM_OUTER_LOOP_54_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_54_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_217_9 = ((ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1);
  assign layer4_out_conc_217_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_217_0 = ((ACCUM_OUTER_LOOP_51_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_51_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_219_9 = ((ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1);
  assign layer4_out_conc_219_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_219_0 = ((ACCUM_OUTER_LOOP_52_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_52_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_221_9 = ((ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1);
  assign layer4_out_conc_221_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_221_0 = ((ACCUM_OUTER_LOOP_49_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_49_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_223_9 = ((ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1);
  assign layer4_out_conc_223_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_223_0 = ((ACCUM_OUTER_LOOP_50_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_50_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_225_9 = ((ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1);
  assign layer4_out_conc_225_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_225_0 = ((ACCUM_OUTER_LOOP_47_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_47_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_227_9 = ((ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1);
  assign layer4_out_conc_227_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_227_0 = ((ACCUM_OUTER_LOOP_48_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_48_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_229_9 = ((ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1);
  assign layer4_out_conc_229_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_229_0 = ((ACCUM_OUTER_LOOP_45_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_45_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_231_9 = ((ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1);
  assign layer4_out_conc_231_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_231_0 = ((ACCUM_OUTER_LOOP_46_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_46_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_233_9 = ((ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1);
  assign layer4_out_conc_233_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_233_0 = ((ACCUM_OUTER_LOOP_43_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_43_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_235_9 = ((ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1);
  assign layer4_out_conc_235_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_235_0 = ((ACCUM_OUTER_LOOP_44_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_44_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_237_9 = ((ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1);
  assign layer4_out_conc_237_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_237_0 = ((ACCUM_OUTER_LOOP_41_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_41_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_239_9 = ((ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1);
  assign layer4_out_conc_239_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_239_0 = ((ACCUM_OUTER_LOOP_42_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_42_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_241_9 = ((ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1);
  assign layer4_out_conc_241_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_241_0 = ((ACCUM_OUTER_LOOP_39_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_39_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_243_9 = ((ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1);
  assign layer4_out_conc_243_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_243_0 = ((ACCUM_OUTER_LOOP_40_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_40_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_245_9 = ((ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1);
  assign layer4_out_conc_245_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_245_0 = ((ACCUM_OUTER_LOOP_37_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_37_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_247_9 = ((ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1);
  assign layer4_out_conc_247_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_247_0 = ((ACCUM_OUTER_LOOP_38_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_38_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_249_9 = ((ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1);
  assign layer4_out_conc_249_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_249_0 = ((ACCUM_OUTER_LOOP_35_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_35_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_251_9 = ((ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1);
  assign layer4_out_conc_251_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_251_0 = ((ACCUM_OUTER_LOOP_36_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_36_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_253_9 = ((ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1);
  assign layer4_out_conc_253_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_253_0 = ((ACCUM_OUTER_LOOP_33_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_33_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_255_9 = ((ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1);
  assign layer4_out_conc_255_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_255_0 = ((ACCUM_OUTER_LOOP_34_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_34_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_257_9 = ((ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1);
  assign layer4_out_conc_257_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_257_0 = ((ACCUM_OUTER_LOOP_31_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_31_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_259_9 = ((ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1);
  assign layer4_out_conc_259_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_259_0 = ((ACCUM_OUTER_LOOP_32_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_32_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_261_9 = ((ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1);
  assign layer4_out_conc_261_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_261_0 = ((ACCUM_OUTER_LOOP_29_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_29_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_263_9 = ((ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1);
  assign layer4_out_conc_263_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_263_0 = ((ACCUM_OUTER_LOOP_30_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_30_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_265_9 = ((ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1);
  assign layer4_out_conc_265_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_265_0 = ((ACCUM_OUTER_LOOP_27_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_27_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_267_9 = ((ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1);
  assign layer4_out_conc_267_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_267_0 = ((ACCUM_OUTER_LOOP_28_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_28_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_269_9 = ((ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1);
  assign layer4_out_conc_269_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_269_0 = ((ACCUM_OUTER_LOOP_25_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_25_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_271_9 = ((ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1);
  assign layer4_out_conc_271_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_271_0 = ((ACCUM_OUTER_LOOP_26_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_26_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_273_9 = ((ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1);
  assign layer4_out_conc_273_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_273_0 = ((ACCUM_OUTER_LOOP_23_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_23_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_275_9 = ((ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1);
  assign layer4_out_conc_275_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_275_0 = ((ACCUM_OUTER_LOOP_24_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_24_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_277_9 = ((ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1);
  assign layer4_out_conc_277_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_277_0 = ((ACCUM_OUTER_LOOP_21_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_21_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_279_9 = ((ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1);
  assign layer4_out_conc_279_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_279_0 = ((ACCUM_OUTER_LOOP_22_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_22_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_281_9 = ((ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1);
  assign layer4_out_conc_281_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_281_0 = ((ACCUM_OUTER_LOOP_19_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_19_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_283_9 = ((ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1);
  assign layer4_out_conc_283_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_283_0 = ((ACCUM_OUTER_LOOP_20_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_20_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_285_9 = ((ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1);
  assign layer4_out_conc_285_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_285_0 = ((ACCUM_OUTER_LOOP_17_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_17_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_287_9 = ((ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1);
  assign layer4_out_conc_287_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_287_0 = ((ACCUM_OUTER_LOOP_18_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_18_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_289_9 = ((ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1);
  assign layer4_out_conc_289_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_289_0 = ((ACCUM_OUTER_LOOP_15_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_15_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_291_9 = ((ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1);
  assign layer4_out_conc_291_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_291_0 = ((ACCUM_OUTER_LOOP_16_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_16_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_293_9 = ((ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1);
  assign layer4_out_conc_293_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_293_0 = ((ACCUM_OUTER_LOOP_13_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_13_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_295_9 = ((ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1);
  assign layer4_out_conc_295_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_295_0 = ((ACCUM_OUTER_LOOP_14_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_14_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_297_9 = ((ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1);
  assign layer4_out_conc_297_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_297_0 = ((ACCUM_OUTER_LOOP_11_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_11_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_299_9 = ((ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1);
  assign layer4_out_conc_299_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_299_0 = ((ACCUM_OUTER_LOOP_12_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_12_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_301_9 = ((ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1);
  assign layer4_out_conc_301_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_301_0 = ((ACCUM_OUTER_LOOP_9_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_9_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_303_9 = ((ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1);
  assign layer4_out_conc_303_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_303_0 = ((ACCUM_OUTER_LOOP_10_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_10_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_305_9 = ((ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1);
  assign layer4_out_conc_305_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_305_0 = ((ACCUM_OUTER_LOOP_7_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_7_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_307_9 = ((ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1);
  assign layer4_out_conc_307_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_307_0 = ((ACCUM_OUTER_LOOP_8_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_8_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_309_9 = ((ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1);
  assign layer4_out_conc_309_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_309_0 = ((ACCUM_OUTER_LOOP_5_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_5_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_311_9 = ((ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1);
  assign layer4_out_conc_311_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_311_0 = ((ACCUM_OUTER_LOOP_6_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_6_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_313_9 = ((ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1);
  assign layer4_out_conc_313_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_313_0 = ((ACCUM_OUTER_LOOP_3_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_3_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_315_9 = ((ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1);
  assign layer4_out_conc_315_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_315_0 = ((ACCUM_OUTER_LOOP_4_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_4_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_317_9 = ((layer2_out_0_sva_1[9]) | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1)
      & nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((layer2_out_0_sva_1[8:1]), 8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1);
  assign layer4_out_conc_317_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_317_0 = ((layer2_out_0_sva_1[0]) | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1)
      & nnet_relu_layer2_t_layer4_t_relu_config4_for_1_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign layer4_out_conc_319_9 = ((ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[9])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  assign nnet_relu_layer2_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl
      = MUX_v_8_2_2((ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[8:1]),
      8'b11111111, nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1);
  assign layer4_out_conc_319_8_1 = MUX_v_8_2_2(8'b00000000, nnet_relu_layer2_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nnet_relu_layer2_t_layer4_t_relu_config4_for_if_or_1_nl,
      nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1);
  assign layer4_out_conc_319_0 = ((ACCUM_OUTER_LOOP_2_ACCUM_INNER_LOOP_14_acc_2_ncse_sva_1[0])
      | nnet_relu_layer2_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1) & nnet_relu_layer2_t_layer4_t_relu_config4_for_2_operator_16_6_true_AC_TRN_AC_WRAP_acc_itm_16_1;
  always @(posedge clk) begin
    if ( rst ) begin
      layer5_out_rsci_idat_15_0 <= 16'b0000000000000000;
      layer5_out_rsci_idat_31_16 <= 16'b0000000000000000;
      layer5_out_rsci_idat_47_32 <= 16'b0000000000000000;
    end
    else begin
      layer5_out_rsci_idat_15_0 <= nl_layer5_out_rsci_idat_15_0[15:0];
      layer5_out_rsci_idat_31_16 <= nl_layer5_out_rsci_idat_31_16[15:0];
      layer5_out_rsci_idat_47_32 <= nl_layer5_out_rsci_idat_47_32[15:0];
    end
  end
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_223_9 , layer4_out_conc_223_8_1 ,
      layer4_out_conc_223_0})) * $signed((w5_rsci_idat[249:245]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_225_9 , layer4_out_conc_225_8_1 ,
      layer4_out_conc_225_0})) * $signed((w5_rsci_idat[234:230]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_227_9 , layer4_out_conc_227_8_1 ,
      layer4_out_conc_227_0})) * $signed((w5_rsci_idat[239:235]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_229_9 , layer4_out_conc_229_8_1 ,
      layer4_out_conc_229_0})) * $signed((w5_rsci_idat[224:220]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_287_9 , layer4_out_conc_287_8_1 ,
      layer4_out_conc_287_0})) * $signed((w5_rsci_idat[89:85]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_289_9 , layer4_out_conc_289_8_1 ,
      layer4_out_conc_289_0})) * $signed((w5_rsci_idat[74:70]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_291_9 , layer4_out_conc_291_8_1 ,
      layer4_out_conc_291_0})) * $signed((w5_rsci_idat[79:75]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_293_9 , layer4_out_conc_293_8_1 ,
      layer4_out_conc_293_0})) * $signed((w5_rsci_idat[64:60]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_295_9 , layer4_out_conc_295_8_1 ,
      layer4_out_conc_295_0})) * $signed((w5_rsci_idat[69:65]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_297_9 , layer4_out_conc_297_8_1 ,
      layer4_out_conc_297_0})) * $signed((w5_rsci_idat[54:50]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_299_9 , layer4_out_conc_299_8_1 ,
      layer4_out_conc_299_0})) * $signed((w5_rsci_idat[59:55]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_301_9 , layer4_out_conc_301_8_1 , layer4_out_conc_301_0}))
      * $signed((w5_rsci_idat[44:40]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_263_9 , layer4_out_conc_263_8_1 ,
      layer4_out_conc_263_0})) * $signed((w5_rsci_idat[149:145]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_265_9 , layer4_out_conc_265_8_1 ,
      layer4_out_conc_265_0})) * $signed((w5_rsci_idat[134:130]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_255_9 , layer4_out_conc_255_8_1 ,
      layer4_out_conc_255_0})) * $signed((w5_rsci_idat[169:165]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_257_9 , layer4_out_conc_257_8_1 ,
      layer4_out_conc_257_0})) * $signed((w5_rsci_idat[154:150]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_259_9 , layer4_out_conc_259_8_1 ,
      layer4_out_conc_259_0})) * $signed((w5_rsci_idat[159:155]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_261_9 , layer4_out_conc_261_8_1 ,
      layer4_out_conc_261_0})) * $signed((w5_rsci_idat[144:140]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_267_9 , layer4_out_conc_267_8_1 ,
      layer4_out_conc_267_0})) * $signed((w5_rsci_idat[139:135]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_269_9 , layer4_out_conc_269_8_1 ,
      layer4_out_conc_269_0})) * $signed((w5_rsci_idat[124:120]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_279_9 , layer4_out_conc_279_8_1 ,
      layer4_out_conc_279_0})) * $signed((w5_rsci_idat[109:105]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_281_9 , layer4_out_conc_281_8_1 ,
      layer4_out_conc_281_0})) * $signed((w5_rsci_idat[94:90]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_271_9 , layer4_out_conc_271_8_1 ,
      layer4_out_conc_271_0})) * $signed((w5_rsci_idat[129:125]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_273_9 , layer4_out_conc_273_8_1 ,
      layer4_out_conc_273_0})) * $signed((w5_rsci_idat[114:110]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_275_9 , layer4_out_conc_275_8_1 ,
      layer4_out_conc_275_0})) * $signed((w5_rsci_idat[119:115]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_277_9 , layer4_out_conc_277_8_1 ,
      layer4_out_conc_277_0})) * $signed((w5_rsci_idat[104:100]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_283_9 , layer4_out_conc_283_8_1 ,
      layer4_out_conc_283_0})) * $signed((w5_rsci_idat[99:95]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_285_9 , layer4_out_conc_285_8_1 ,
      layer4_out_conc_285_0})) * $signed((w5_rsci_idat[84:80]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_0}))
      * $signed((w5_rsci_idat[329:325]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_193_9 , layer4_out_conc_193_8_1 ,
      layer4_out_conc_193_0})) * $signed((w5_rsci_idat[314:310]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_195_9 , layer4_out_conc_195_8_1 ,
      layer4_out_conc_195_0})) * $signed((w5_rsci_idat[319:315]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_197_9 , layer4_out_conc_197_8_1 ,
      layer4_out_conc_197_0})) * $signed((w5_rsci_idat[304:300]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_199_9 , layer4_out_conc_199_8_1 ,
      layer4_out_conc_199_0})) * $signed((w5_rsci_idat[309:305]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_201_9 , layer4_out_conc_201_8_1 ,
      layer4_out_conc_201_0})) * $signed((w5_rsci_idat[294:290]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_203_9 , layer4_out_conc_203_8_1 ,
      layer4_out_conc_203_0})) * $signed((w5_rsci_idat[299:295]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_205_9 , layer4_out_conc_205_8_1 ,
      layer4_out_conc_205_0})) * $signed((w5_rsci_idat[284:280]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_215_9 , layer4_out_conc_215_8_1 ,
      layer4_out_conc_215_0})) * $signed((w5_rsci_idat[269:265]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_217_9 , layer4_out_conc_217_8_1 ,
      layer4_out_conc_217_0})) * $signed((w5_rsci_idat[254:250]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_219_9 , layer4_out_conc_219_8_1 ,
      layer4_out_conc_219_0})) * $signed((w5_rsci_idat[259:255]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_221_9 , layer4_out_conc_221_8_1 ,
      layer4_out_conc_221_0})) * $signed((w5_rsci_idat[244:240]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_207_9 , layer4_out_conc_207_8_1 ,
      layer4_out_conc_207_0})) * $signed((w5_rsci_idat[289:285]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_209_9 , layer4_out_conc_209_8_1 ,
      layer4_out_conc_209_0})) * $signed((w5_rsci_idat[274:270]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_211_9 , layer4_out_conc_211_8_1 ,
      layer4_out_conc_211_0})) * $signed((w5_rsci_idat[279:275]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_213_9 , layer4_out_conc_213_8_1 ,
      layer4_out_conc_213_0})) * $signed((w5_rsci_idat[264:260]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_231_9 , layer4_out_conc_231_8_1 ,
      layer4_out_conc_231_0})) * $signed((w5_rsci_idat[229:225]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_233_9 , layer4_out_conc_233_8_1 ,
      layer4_out_conc_233_0})) * $signed((w5_rsci_idat[214:210]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_235_9 , layer4_out_conc_235_8_1 ,
      layer4_out_conc_235_0})) * $signed((w5_rsci_idat[219:215]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_237_9 , layer4_out_conc_237_8_1 ,
      layer4_out_conc_237_0})) * $signed((w5_rsci_idat[204:200]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_247_9 , layer4_out_conc_247_8_1 ,
      layer4_out_conc_247_0})) * $signed((w5_rsci_idat[189:185]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_249_9 , layer4_out_conc_249_8_1 ,
      layer4_out_conc_249_0})) * $signed((w5_rsci_idat[174:170]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_251_9 , layer4_out_conc_251_8_1 ,
      layer4_out_conc_251_0})) * $signed((w5_rsci_idat[179:175]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_253_9 , layer4_out_conc_253_8_1 ,
      layer4_out_conc_253_0})) * $signed((w5_rsci_idat[164:160]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_239_9 , layer4_out_conc_239_8_1 ,
      layer4_out_conc_239_0})) * $signed((w5_rsci_idat[209:205]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_241_9 , layer4_out_conc_241_8_1 ,
      layer4_out_conc_241_0})) * $signed((w5_rsci_idat[194:190]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_243_9 , layer4_out_conc_243_8_1 ,
      layer4_out_conc_243_0})) * $signed((w5_rsci_idat[199:195]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_245_9 , layer4_out_conc_245_8_1 ,
      layer4_out_conc_245_0})) * $signed((w5_rsci_idat[184:180]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_311_9 , layer4_out_conc_311_8_1 , layer4_out_conc_311_0}))
      * $signed((w5_rsci_idat[29:25]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_313_9 , layer4_out_conc_313_8_1 , layer4_out_conc_313_0}))
      * $signed((w5_rsci_idat[14:10]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_315_9 , layer4_out_conc_315_8_1 , layer4_out_conc_315_0}))
      * $signed((w5_rsci_idat[19:15]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_317_9 , layer4_out_conc_317_8_1 , layer4_out_conc_317_0}))
      * $signed((w5_rsci_idat[4:0]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_303_9 , layer4_out_conc_303_8_1 ,
      layer4_out_conc_303_0})) * $signed((w5_rsci_idat[49:45]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_305_9 , layer4_out_conc_305_8_1 , layer4_out_conc_305_0}))
      * $signed((w5_rsci_idat[34:30]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_307_9 , layer4_out_conc_307_8_1 , layer4_out_conc_307_0}))
      * $signed((w5_rsci_idat[39:35]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_309_9 , layer4_out_conc_309_8_1 , layer4_out_conc_309_0}))
      * $signed((w5_rsci_idat[24:20]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_393_nl = conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl));
  assign ACCUM_INNER_LOOP_1_acc_393_nl = nl_ACCUM_INNER_LOOP_1_acc_393_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_0}))
      * $signed((w5_rsci_idat[629:625]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_0}))
      * $signed((w5_rsci_idat[614:610]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_0}))
      * $signed((w5_rsci_idat[589:585]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_0}))
      * $signed((w5_rsci_idat[574:570]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_0}))
      * $signed((w5_rsci_idat[609:605]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_0}))
      * $signed((w5_rsci_idat[594:590]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_0}))
      * $signed((w5_rsci_idat[509:505]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_0}))
      * $signed((w5_rsci_idat[494:490]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_0}))
      * $signed((w5_rsci_idat[529:525]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_0}))
      * $signed((w5_rsci_idat[514:510]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_0}))
      * $signed((w5_rsci_idat[519:515]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_0}))
      * $signed((w5_rsci_idat[504:500]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_0}))
      * $signed((w5_rsci_idat[569:565]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_0}))
      * $signed((w5_rsci_idat[554:550]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_0}))
      * $signed((w5_rsci_idat[559:555]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_0}))
      * $signed((w5_rsci_idat[544:540]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_0}))
      * $signed((w5_rsci_idat[549:545]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_0}))
      * $signed((w5_rsci_idat[534:530]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_0}))
      * $signed((w5_rsci_idat[539:535]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_0}))
      * $signed((w5_rsci_idat[524:520]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_396_nl = conv_s2s_5_6(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1[10:6])
      + conv_s2s_5_6(b5_rsci_idat[4:0]);
  assign ACCUM_INNER_LOOP_1_acc_396_nl = nl_ACCUM_INNER_LOOP_1_acc_396_nl[5:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_0}))
      * $signed((w5_rsci_idat[634:630]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_0}))
      * $signed((w5_rsci_idat[639:635]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_0}))
      * $signed((w5_rsci_idat[624:620]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_0}))
      * $signed((w5_rsci_idat[619:615]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_0}))
      * $signed((w5_rsci_idat[604:600]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_0}))
      * $signed((w5_rsci_idat[599:595]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_0}))
      * $signed((w5_rsci_idat[584:580]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_0}))
      * $signed((w5_rsci_idat[579:575]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_0}))
      * $signed((w5_rsci_idat[564:560]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_0}))
      * $signed((w5_rsci_idat[499:495]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_0}))
      * $signed((w5_rsci_idat[484:480]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_392_nl = conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_12_16({ACCUM_INNER_LOOP_1_acc_396_nl , (ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1[5:0])})
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl));
  assign ACCUM_INNER_LOOP_1_acc_392_nl = nl_ACCUM_INNER_LOOP_1_acc_392_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_0}))
      * $signed((w5_rsci_idat[469:465]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_0}))
      * $signed((w5_rsci_idat[454:450]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_0}))
      * $signed((w5_rsci_idat[489:485]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_0}))
      * $signed((w5_rsci_idat[474:470]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_0}))
      * $signed((w5_rsci_idat[429:425]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_0}))
      * $signed((w5_rsci_idat[414:410]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_0}))
      * $signed((w5_rsci_idat[449:445]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_0}))
      * $signed((w5_rsci_idat[434:430]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_0}))
      * $signed((w5_rsci_idat[439:435]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_0}))
      * $signed((w5_rsci_idat[424:420]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_0}))
      * $signed((w5_rsci_idat[409:405]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_0}))
      * $signed((w5_rsci_idat[394:390]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_0}))
      * $signed((w5_rsci_idat[399:395]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_0}))
      * $signed((w5_rsci_idat[384:380]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_0}))
      * $signed((w5_rsci_idat[389:385]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_0}))
      * $signed((w5_rsci_idat[374:370]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_0}))
      * $signed((w5_rsci_idat[379:375]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_0}))
      * $signed((w5_rsci_idat[364:360]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_0}))
      * $signed((w5_rsci_idat[349:345]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_0}))
      * $signed((w5_rsci_idat[334:330]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_0}))
      * $signed((w5_rsci_idat[339:335]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_0}))
      * $signed((w5_rsci_idat[324:320]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_0}))
      * $signed((w5_rsci_idat[369:365]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_0}))
      * $signed((w5_rsci_idat[354:350]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_0}))
      * $signed((w5_rsci_idat[359:355]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_0}))
      * $signed((w5_rsci_idat[344:340]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_0}))
      * $signed((w5_rsci_idat[479:475]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_0}))
      * $signed((w5_rsci_idat[464:460]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_0}))
      * $signed((w5_rsci_idat[459:455]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_0}))
      * $signed((w5_rsci_idat[444:440]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_0}))
      * $signed((w5_rsci_idat[419:415]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_0}))
      * $signed((w5_rsci_idat[404:400]));
  assign ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_layer5_out_rsci_idat_15_0  = ACCUM_INNER_LOOP_1_acc_393_nl + ACCUM_INNER_LOOP_1_acc_392_nl
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_1_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl));
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_223_9 , layer4_out_conc_223_8_1 ,
      layer4_out_conc_223_0})) * $signed((w5_rsci_idat[889:885]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_225_9 , layer4_out_conc_225_8_1 ,
      layer4_out_conc_225_0})) * $signed((w5_rsci_idat[874:870]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_227_9 , layer4_out_conc_227_8_1 ,
      layer4_out_conc_227_0})) * $signed((w5_rsci_idat[879:875]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_229_9 , layer4_out_conc_229_8_1 ,
      layer4_out_conc_229_0})) * $signed((w5_rsci_idat[864:860]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_287_9 , layer4_out_conc_287_8_1 ,
      layer4_out_conc_287_0})) * $signed((w5_rsci_idat[729:725]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_289_9 , layer4_out_conc_289_8_1 ,
      layer4_out_conc_289_0})) * $signed((w5_rsci_idat[714:710]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_291_9 , layer4_out_conc_291_8_1 ,
      layer4_out_conc_291_0})) * $signed((w5_rsci_idat[719:715]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_293_9 , layer4_out_conc_293_8_1 ,
      layer4_out_conc_293_0})) * $signed((w5_rsci_idat[704:700]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_295_9 , layer4_out_conc_295_8_1 ,
      layer4_out_conc_295_0})) * $signed((w5_rsci_idat[709:705]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_297_9 , layer4_out_conc_297_8_1 ,
      layer4_out_conc_297_0})) * $signed((w5_rsci_idat[694:690]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_299_9 , layer4_out_conc_299_8_1 ,
      layer4_out_conc_299_0})) * $signed((w5_rsci_idat[699:695]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_301_9 , layer4_out_conc_301_8_1 , layer4_out_conc_301_0}))
      * $signed((w5_rsci_idat[684:680]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_263_9 , layer4_out_conc_263_8_1 ,
      layer4_out_conc_263_0})) * $signed((w5_rsci_idat[789:785]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_265_9 , layer4_out_conc_265_8_1 ,
      layer4_out_conc_265_0})) * $signed((w5_rsci_idat[774:770]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_255_9 , layer4_out_conc_255_8_1 ,
      layer4_out_conc_255_0})) * $signed((w5_rsci_idat[809:805]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_257_9 , layer4_out_conc_257_8_1 ,
      layer4_out_conc_257_0})) * $signed((w5_rsci_idat[794:790]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_259_9 , layer4_out_conc_259_8_1 ,
      layer4_out_conc_259_0})) * $signed((w5_rsci_idat[799:795]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_261_9 , layer4_out_conc_261_8_1 ,
      layer4_out_conc_261_0})) * $signed((w5_rsci_idat[784:780]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_267_9 , layer4_out_conc_267_8_1 ,
      layer4_out_conc_267_0})) * $signed((w5_rsci_idat[779:775]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_269_9 , layer4_out_conc_269_8_1 ,
      layer4_out_conc_269_0})) * $signed((w5_rsci_idat[764:760]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_279_9 , layer4_out_conc_279_8_1 ,
      layer4_out_conc_279_0})) * $signed((w5_rsci_idat[749:745]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_281_9 , layer4_out_conc_281_8_1 ,
      layer4_out_conc_281_0})) * $signed((w5_rsci_idat[734:730]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_271_9 , layer4_out_conc_271_8_1 ,
      layer4_out_conc_271_0})) * $signed((w5_rsci_idat[769:765]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_273_9 , layer4_out_conc_273_8_1 ,
      layer4_out_conc_273_0})) * $signed((w5_rsci_idat[754:750]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_275_9 , layer4_out_conc_275_8_1 ,
      layer4_out_conc_275_0})) * $signed((w5_rsci_idat[759:755]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_277_9 , layer4_out_conc_277_8_1 ,
      layer4_out_conc_277_0})) * $signed((w5_rsci_idat[744:740]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_283_9 , layer4_out_conc_283_8_1 ,
      layer4_out_conc_283_0})) * $signed((w5_rsci_idat[739:735]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_285_9 , layer4_out_conc_285_8_1 ,
      layer4_out_conc_285_0})) * $signed((w5_rsci_idat[724:720]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_0}))
      * $signed((w5_rsci_idat[969:965]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_193_9 , layer4_out_conc_193_8_1 ,
      layer4_out_conc_193_0})) * $signed((w5_rsci_idat[954:950]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_195_9 , layer4_out_conc_195_8_1 ,
      layer4_out_conc_195_0})) * $signed((w5_rsci_idat[959:955]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_197_9 , layer4_out_conc_197_8_1 ,
      layer4_out_conc_197_0})) * $signed((w5_rsci_idat[944:940]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_199_9 , layer4_out_conc_199_8_1 ,
      layer4_out_conc_199_0})) * $signed((w5_rsci_idat[949:945]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_201_9 , layer4_out_conc_201_8_1 ,
      layer4_out_conc_201_0})) * $signed((w5_rsci_idat[934:930]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_203_9 , layer4_out_conc_203_8_1 ,
      layer4_out_conc_203_0})) * $signed((w5_rsci_idat[939:935]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_205_9 , layer4_out_conc_205_8_1 ,
      layer4_out_conc_205_0})) * $signed((w5_rsci_idat[924:920]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_215_9 , layer4_out_conc_215_8_1 ,
      layer4_out_conc_215_0})) * $signed((w5_rsci_idat[909:905]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_217_9 , layer4_out_conc_217_8_1 ,
      layer4_out_conc_217_0})) * $signed((w5_rsci_idat[894:890]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_219_9 , layer4_out_conc_219_8_1 ,
      layer4_out_conc_219_0})) * $signed((w5_rsci_idat[899:895]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_221_9 , layer4_out_conc_221_8_1 ,
      layer4_out_conc_221_0})) * $signed((w5_rsci_idat[884:880]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_207_9 , layer4_out_conc_207_8_1 ,
      layer4_out_conc_207_0})) * $signed((w5_rsci_idat[929:925]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_209_9 , layer4_out_conc_209_8_1 ,
      layer4_out_conc_209_0})) * $signed((w5_rsci_idat[914:910]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_211_9 , layer4_out_conc_211_8_1 ,
      layer4_out_conc_211_0})) * $signed((w5_rsci_idat[919:915]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_213_9 , layer4_out_conc_213_8_1 ,
      layer4_out_conc_213_0})) * $signed((w5_rsci_idat[904:900]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_231_9 , layer4_out_conc_231_8_1 ,
      layer4_out_conc_231_0})) * $signed((w5_rsci_idat[869:865]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_233_9 , layer4_out_conc_233_8_1 ,
      layer4_out_conc_233_0})) * $signed((w5_rsci_idat[854:850]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_235_9 , layer4_out_conc_235_8_1 ,
      layer4_out_conc_235_0})) * $signed((w5_rsci_idat[859:855]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_237_9 , layer4_out_conc_237_8_1 ,
      layer4_out_conc_237_0})) * $signed((w5_rsci_idat[844:840]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_247_9 , layer4_out_conc_247_8_1 ,
      layer4_out_conc_247_0})) * $signed((w5_rsci_idat[829:825]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_249_9 , layer4_out_conc_249_8_1 ,
      layer4_out_conc_249_0})) * $signed((w5_rsci_idat[814:810]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_251_9 , layer4_out_conc_251_8_1 ,
      layer4_out_conc_251_0})) * $signed((w5_rsci_idat[819:815]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_253_9 , layer4_out_conc_253_8_1 ,
      layer4_out_conc_253_0})) * $signed((w5_rsci_idat[804:800]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_239_9 , layer4_out_conc_239_8_1 ,
      layer4_out_conc_239_0})) * $signed((w5_rsci_idat[849:845]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_241_9 , layer4_out_conc_241_8_1 ,
      layer4_out_conc_241_0})) * $signed((w5_rsci_idat[834:830]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_243_9 , layer4_out_conc_243_8_1 ,
      layer4_out_conc_243_0})) * $signed((w5_rsci_idat[839:835]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_245_9 , layer4_out_conc_245_8_1 ,
      layer4_out_conc_245_0})) * $signed((w5_rsci_idat[824:820]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_311_9 , layer4_out_conc_311_8_1 , layer4_out_conc_311_0}))
      * $signed((w5_rsci_idat[669:665]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_313_9 , layer4_out_conc_313_8_1 , layer4_out_conc_313_0}))
      * $signed((w5_rsci_idat[654:650]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_315_9 , layer4_out_conc_315_8_1 , layer4_out_conc_315_0}))
      * $signed((w5_rsci_idat[659:655]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_317_9 , layer4_out_conc_317_8_1 , layer4_out_conc_317_0}))
      * $signed((w5_rsci_idat[644:640]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_303_9 , layer4_out_conc_303_8_1 ,
      layer4_out_conc_303_0})) * $signed((w5_rsci_idat[689:685]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_305_9 , layer4_out_conc_305_8_1 , layer4_out_conc_305_0}))
      * $signed((w5_rsci_idat[674:670]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_307_9 , layer4_out_conc_307_8_1 , layer4_out_conc_307_0}))
      * $signed((w5_rsci_idat[679:675]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_309_9 , layer4_out_conc_309_8_1 , layer4_out_conc_309_0}))
      * $signed((w5_rsci_idat[664:660]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_266_nl = conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl));
  assign ACCUM_INNER_LOOP_1_acc_266_nl = nl_ACCUM_INNER_LOOP_1_acc_266_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_0}))
      * $signed((w5_rsci_idat[1269:1265]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_0}))
      * $signed((w5_rsci_idat[1254:1250]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_0}))
      * $signed((w5_rsci_idat[1229:1225]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_0}))
      * $signed((w5_rsci_idat[1214:1210]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_0}))
      * $signed((w5_rsci_idat[1249:1245]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_0}))
      * $signed((w5_rsci_idat[1234:1230]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_0}))
      * $signed((w5_rsci_idat[1149:1145]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_0}))
      * $signed((w5_rsci_idat[1134:1130]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_0}))
      * $signed((w5_rsci_idat[1169:1165]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_0}))
      * $signed((w5_rsci_idat[1154:1150]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_0}))
      * $signed((w5_rsci_idat[1159:1155]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_0}))
      * $signed((w5_rsci_idat[1144:1140]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_0}))
      * $signed((w5_rsci_idat[1209:1205]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_0}))
      * $signed((w5_rsci_idat[1194:1190]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_0}))
      * $signed((w5_rsci_idat[1199:1195]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_0}))
      * $signed((w5_rsci_idat[1184:1180]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_0}))
      * $signed((w5_rsci_idat[1189:1185]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_0}))
      * $signed((w5_rsci_idat[1174:1170]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_0}))
      * $signed((w5_rsci_idat[1179:1175]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_0}))
      * $signed((w5_rsci_idat[1164:1160]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_395_nl = conv_s2s_5_6(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1[10:6])
      + conv_s2s_5_6(b5_rsci_idat[9:5]);
  assign ACCUM_INNER_LOOP_1_acc_395_nl = nl_ACCUM_INNER_LOOP_1_acc_395_nl[5:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_0}))
      * $signed((w5_rsci_idat[1274:1270]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_0}))
      * $signed((w5_rsci_idat[1279:1275]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_0}))
      * $signed((w5_rsci_idat[1264:1260]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_0}))
      * $signed((w5_rsci_idat[1259:1255]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_0}))
      * $signed((w5_rsci_idat[1244:1240]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_0}))
      * $signed((w5_rsci_idat[1239:1235]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_0}))
      * $signed((w5_rsci_idat[1224:1220]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_0}))
      * $signed((w5_rsci_idat[1219:1215]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_0}))
      * $signed((w5_rsci_idat[1204:1200]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_0}))
      * $signed((w5_rsci_idat[1139:1135]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_0}))
      * $signed((w5_rsci_idat[1124:1120]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_265_nl = conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_12_16({ACCUM_INNER_LOOP_1_acc_395_nl , (ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1[5:0])})
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl));
  assign ACCUM_INNER_LOOP_1_acc_265_nl = nl_ACCUM_INNER_LOOP_1_acc_265_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_0}))
      * $signed((w5_rsci_idat[1109:1105]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_0}))
      * $signed((w5_rsci_idat[1094:1090]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_0}))
      * $signed((w5_rsci_idat[1129:1125]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_0}))
      * $signed((w5_rsci_idat[1114:1110]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_0}))
      * $signed((w5_rsci_idat[1069:1065]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_0}))
      * $signed((w5_rsci_idat[1054:1050]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_0}))
      * $signed((w5_rsci_idat[1089:1085]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_0}))
      * $signed((w5_rsci_idat[1074:1070]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_0}))
      * $signed((w5_rsci_idat[1079:1075]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_0}))
      * $signed((w5_rsci_idat[1064:1060]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_0}))
      * $signed((w5_rsci_idat[1049:1045]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_0}))
      * $signed((w5_rsci_idat[1034:1030]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_0}))
      * $signed((w5_rsci_idat[1039:1035]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_0}))
      * $signed((w5_rsci_idat[1024:1020]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_0}))
      * $signed((w5_rsci_idat[1029:1025]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_0}))
      * $signed((w5_rsci_idat[1014:1010]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_0}))
      * $signed((w5_rsci_idat[1019:1015]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_0}))
      * $signed((w5_rsci_idat[1004:1000]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_0}))
      * $signed((w5_rsci_idat[989:985]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_0}))
      * $signed((w5_rsci_idat[974:970]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_0}))
      * $signed((w5_rsci_idat[979:975]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_0}))
      * $signed((w5_rsci_idat[964:960]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_0}))
      * $signed((w5_rsci_idat[1009:1005]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_0}))
      * $signed((w5_rsci_idat[994:990]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_0}))
      * $signed((w5_rsci_idat[999:995]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_0}))
      * $signed((w5_rsci_idat[984:980]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_0}))
      * $signed((w5_rsci_idat[1119:1115]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_0}))
      * $signed((w5_rsci_idat[1104:1100]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_0}))
      * $signed((w5_rsci_idat[1099:1095]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_0}))
      * $signed((w5_rsci_idat[1084:1080]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_0}))
      * $signed((w5_rsci_idat[1059:1055]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_0}))
      * $signed((w5_rsci_idat[1044:1040]));
  assign ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_layer5_out_rsci_idat_31_16  = ACCUM_INNER_LOOP_1_acc_266_nl + ACCUM_INNER_LOOP_1_acc_265_nl
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_2_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl));
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_223_9 , layer4_out_conc_223_8_1 ,
      layer4_out_conc_223_0})) * $signed((w5_rsci_idat[1529:1525]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_225_9 , layer4_out_conc_225_8_1 ,
      layer4_out_conc_225_0})) * $signed((w5_rsci_idat[1514:1510]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_227_9 , layer4_out_conc_227_8_1 ,
      layer4_out_conc_227_0})) * $signed((w5_rsci_idat[1519:1515]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_229_9 , layer4_out_conc_229_8_1 ,
      layer4_out_conc_229_0})) * $signed((w5_rsci_idat[1504:1500]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_287_9 , layer4_out_conc_287_8_1 ,
      layer4_out_conc_287_0})) * $signed((w5_rsci_idat[1369:1365]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_289_9 , layer4_out_conc_289_8_1 ,
      layer4_out_conc_289_0})) * $signed((w5_rsci_idat[1354:1350]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_291_9 , layer4_out_conc_291_8_1 ,
      layer4_out_conc_291_0})) * $signed((w5_rsci_idat[1359:1355]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_293_9 , layer4_out_conc_293_8_1 ,
      layer4_out_conc_293_0})) * $signed((w5_rsci_idat[1344:1340]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_295_9 , layer4_out_conc_295_8_1 ,
      layer4_out_conc_295_0})) * $signed((w5_rsci_idat[1349:1345]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_297_9 , layer4_out_conc_297_8_1 ,
      layer4_out_conc_297_0})) * $signed((w5_rsci_idat[1334:1330]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_299_9 , layer4_out_conc_299_8_1 ,
      layer4_out_conc_299_0})) * $signed((w5_rsci_idat[1339:1335]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_301_9 , layer4_out_conc_301_8_1 , layer4_out_conc_301_0}))
      * $signed((w5_rsci_idat[1324:1320]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_263_9 , layer4_out_conc_263_8_1 ,
      layer4_out_conc_263_0})) * $signed((w5_rsci_idat[1429:1425]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_265_9 , layer4_out_conc_265_8_1 ,
      layer4_out_conc_265_0})) * $signed((w5_rsci_idat[1414:1410]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_255_9 , layer4_out_conc_255_8_1 ,
      layer4_out_conc_255_0})) * $signed((w5_rsci_idat[1449:1445]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_257_9 , layer4_out_conc_257_8_1 ,
      layer4_out_conc_257_0})) * $signed((w5_rsci_idat[1434:1430]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_259_9 , layer4_out_conc_259_8_1 ,
      layer4_out_conc_259_0})) * $signed((w5_rsci_idat[1439:1435]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_261_9 , layer4_out_conc_261_8_1 ,
      layer4_out_conc_261_0})) * $signed((w5_rsci_idat[1424:1420]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_267_9 , layer4_out_conc_267_8_1 ,
      layer4_out_conc_267_0})) * $signed((w5_rsci_idat[1419:1415]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_269_9 , layer4_out_conc_269_8_1 ,
      layer4_out_conc_269_0})) * $signed((w5_rsci_idat[1404:1400]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_279_9 , layer4_out_conc_279_8_1 ,
      layer4_out_conc_279_0})) * $signed((w5_rsci_idat[1389:1385]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_281_9 , layer4_out_conc_281_8_1 ,
      layer4_out_conc_281_0})) * $signed((w5_rsci_idat[1374:1370]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_271_9 , layer4_out_conc_271_8_1 ,
      layer4_out_conc_271_0})) * $signed((w5_rsci_idat[1409:1405]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_273_9 , layer4_out_conc_273_8_1 ,
      layer4_out_conc_273_0})) * $signed((w5_rsci_idat[1394:1390]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_275_9 , layer4_out_conc_275_8_1 ,
      layer4_out_conc_275_0})) * $signed((w5_rsci_idat[1399:1395]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_277_9 , layer4_out_conc_277_8_1 ,
      layer4_out_conc_277_0})) * $signed((w5_rsci_idat[1384:1380]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_283_9 , layer4_out_conc_283_8_1 ,
      layer4_out_conc_283_0})) * $signed((w5_rsci_idat[1379:1375]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_285_9 , layer4_out_conc_285_8_1 ,
      layer4_out_conc_285_0})) * $signed((w5_rsci_idat[1364:1360]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_384_0}))
      * $signed((w5_rsci_idat[1609:1605]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_193_9 , layer4_out_conc_193_8_1 ,
      layer4_out_conc_193_0})) * $signed((w5_rsci_idat[1594:1590]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_195_9 , layer4_out_conc_195_8_1 ,
      layer4_out_conc_195_0})) * $signed((w5_rsci_idat[1599:1595]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_197_9 , layer4_out_conc_197_8_1 ,
      layer4_out_conc_197_0})) * $signed((w5_rsci_idat[1584:1580]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_199_9 , layer4_out_conc_199_8_1 ,
      layer4_out_conc_199_0})) * $signed((w5_rsci_idat[1589:1585]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_201_9 , layer4_out_conc_201_8_1 ,
      layer4_out_conc_201_0})) * $signed((w5_rsci_idat[1574:1570]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_203_9 , layer4_out_conc_203_8_1 ,
      layer4_out_conc_203_0})) * $signed((w5_rsci_idat[1579:1575]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_205_9 , layer4_out_conc_205_8_1 ,
      layer4_out_conc_205_0})) * $signed((w5_rsci_idat[1564:1560]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_215_9 , layer4_out_conc_215_8_1 ,
      layer4_out_conc_215_0})) * $signed((w5_rsci_idat[1549:1545]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_217_9 , layer4_out_conc_217_8_1 ,
      layer4_out_conc_217_0})) * $signed((w5_rsci_idat[1534:1530]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_219_9 , layer4_out_conc_219_8_1 ,
      layer4_out_conc_219_0})) * $signed((w5_rsci_idat[1539:1535]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_221_9 , layer4_out_conc_221_8_1 ,
      layer4_out_conc_221_0})) * $signed((w5_rsci_idat[1524:1520]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_207_9 , layer4_out_conc_207_8_1 ,
      layer4_out_conc_207_0})) * $signed((w5_rsci_idat[1569:1565]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_209_9 , layer4_out_conc_209_8_1 ,
      layer4_out_conc_209_0})) * $signed((w5_rsci_idat[1554:1550]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_211_9 , layer4_out_conc_211_8_1 ,
      layer4_out_conc_211_0})) * $signed((w5_rsci_idat[1559:1555]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_213_9 , layer4_out_conc_213_8_1 ,
      layer4_out_conc_213_0})) * $signed((w5_rsci_idat[1544:1540]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_231_9 , layer4_out_conc_231_8_1 ,
      layer4_out_conc_231_0})) * $signed((w5_rsci_idat[1509:1505]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_233_9 , layer4_out_conc_233_8_1 ,
      layer4_out_conc_233_0})) * $signed((w5_rsci_idat[1494:1490]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_235_9 , layer4_out_conc_235_8_1 ,
      layer4_out_conc_235_0})) * $signed((w5_rsci_idat[1499:1495]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_237_9 , layer4_out_conc_237_8_1 ,
      layer4_out_conc_237_0})) * $signed((w5_rsci_idat[1484:1480]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_247_9 , layer4_out_conc_247_8_1 ,
      layer4_out_conc_247_0})) * $signed((w5_rsci_idat[1469:1465]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_249_9 , layer4_out_conc_249_8_1 ,
      layer4_out_conc_249_0})) * $signed((w5_rsci_idat[1454:1450]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_251_9 , layer4_out_conc_251_8_1 ,
      layer4_out_conc_251_0})) * $signed((w5_rsci_idat[1459:1455]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_253_9 , layer4_out_conc_253_8_1 ,
      layer4_out_conc_253_0})) * $signed((w5_rsci_idat[1444:1440]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_239_9 , layer4_out_conc_239_8_1 ,
      layer4_out_conc_239_0})) * $signed((w5_rsci_idat[1489:1485]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_241_9 , layer4_out_conc_241_8_1 ,
      layer4_out_conc_241_0})) * $signed((w5_rsci_idat[1474:1470]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_243_9 , layer4_out_conc_243_8_1 ,
      layer4_out_conc_243_0})) * $signed((w5_rsci_idat[1479:1475]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_245_9 , layer4_out_conc_245_8_1 ,
      layer4_out_conc_245_0})) * $signed((w5_rsci_idat[1464:1460]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_311_9 , layer4_out_conc_311_8_1 , layer4_out_conc_311_0}))
      * $signed((w5_rsci_idat[1309:1305]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_313_9 , layer4_out_conc_313_8_1 , layer4_out_conc_313_0}))
      * $signed((w5_rsci_idat[1294:1290]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_315_9 , layer4_out_conc_315_8_1 , layer4_out_conc_315_0}))
      * $signed((w5_rsci_idat[1299:1295]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_317_9 , layer4_out_conc_317_8_1 , layer4_out_conc_317_0}))
      * $signed((w5_rsci_idat[1284:1280]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_303_9 , layer4_out_conc_303_8_1 ,
      layer4_out_conc_303_0})) * $signed((w5_rsci_idat[1329:1325]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_305_9 , layer4_out_conc_305_8_1 , layer4_out_conc_305_0}))
      * $signed((w5_rsci_idat[1314:1310]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_307_9 , layer4_out_conc_307_8_1 , layer4_out_conc_307_0}))
      * $signed((w5_rsci_idat[1319:1315]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl =
      $signed(conv_u2s_10_11({layer4_out_conc_309_9 , layer4_out_conc_309_8_1 , layer4_out_conc_309_0}))
      * $signed((w5_rsci_idat[1304:1300]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_139_nl = conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_50_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_47_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_48_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_45_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_18_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_15_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_16_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_13_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_14_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_11_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_12_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_9_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_30_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_27_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_34_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_31_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_32_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_29_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_28_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_25_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_22_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_19_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_26_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_23_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_24_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_21_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_20_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_17_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_66_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_63_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_64_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_61_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_62_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_59_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_60_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_57_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_54_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_51_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_52_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_49_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_58_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_55_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_56_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_53_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_46_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_43_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_44_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_41_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_38_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_35_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_36_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_33_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_42_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_39_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_40_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_37_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_6_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_3_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_4_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_1_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_10_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_7_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_8_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_5_ACCUM_INNER_LOOP_1_mul_nl));
  assign ACCUM_INNER_LOOP_1_acc_139_nl = nl_ACCUM_INNER_LOOP_1_acc_139_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_264_0}))
      * $signed((w5_rsci_idat[1909:1905]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_266_0}))
      * $signed((w5_rsci_idat[1894:1890]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_280_0}))
      * $signed((w5_rsci_idat[1869:1865]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_282_0}))
      * $signed((w5_rsci_idat[1854:1850]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_272_0}))
      * $signed((w5_rsci_idat[1889:1885]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_274_0}))
      * $signed((w5_rsci_idat[1874:1870]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_312_0}))
      * $signed((w5_rsci_idat[1789:1785]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_314_0}))
      * $signed((w5_rsci_idat[1774:1770]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_304_0}))
      * $signed((w5_rsci_idat[1809:1805]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_306_0}))
      * $signed((w5_rsci_idat[1794:1790]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_308_0}))
      * $signed((w5_rsci_idat[1799:1795]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_310_0}))
      * $signed((w5_rsci_idat[1784:1780]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_288_0}))
      * $signed((w5_rsci_idat[1849:1845]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_290_0}))
      * $signed((w5_rsci_idat[1834:1830]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_292_0}))
      * $signed((w5_rsci_idat[1839:1835]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_294_0}))
      * $signed((w5_rsci_idat[1824:1820]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_296_0}))
      * $signed((w5_rsci_idat[1829:1825]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_298_0}))
      * $signed((w5_rsci_idat[1814:1810]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_300_0}))
      * $signed((w5_rsci_idat[1819:1815]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_302_0}))
      * $signed((w5_rsci_idat[1804:1800]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_397_nl = conv_s2s_5_6(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1[10:6])
      + conv_s2s_5_6(b5_rsci_idat[14:10]);
  assign ACCUM_INNER_LOOP_1_acc_397_nl = nl_ACCUM_INNER_LOOP_1_acc_397_nl[5:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_258_0}))
      * $signed((w5_rsci_idat[1914:1910]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_260_0}))
      * $signed((w5_rsci_idat[1919:1915]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_262_0}))
      * $signed((w5_rsci_idat[1904:1900]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_268_0}))
      * $signed((w5_rsci_idat[1899:1895]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_270_0}))
      * $signed((w5_rsci_idat[1884:1880]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_276_0}))
      * $signed((w5_rsci_idat[1879:1875]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_278_0}))
      * $signed((w5_rsci_idat[1864:1860]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_284_0}))
      * $signed((w5_rsci_idat[1859:1855]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_286_0}))
      * $signed((w5_rsci_idat[1844:1840]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_316_0}))
      * $signed((w5_rsci_idat[1779:1775]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl =
      nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_318_0}))
      * $signed((w5_rsci_idat[1764:1760]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_INNER_LOOP_1_acc_140_nl = conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_126_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_123_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_118_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_115_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_122_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_119_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_102_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_99_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_106_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_103_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_104_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_101_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_114_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_111_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_112_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_109_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_110_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_107_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_108_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_105_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_12_16({ACCUM_INNER_LOOP_1_acc_397_nl , (ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_2_ACCUM_INNER_LOOP_1_mul_itm_14_4_1[5:0])})
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_127_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_128_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_125_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_124_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_121_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_120_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_117_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_116_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_113_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_100_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_97_ACCUM_INNER_LOOP_1_mul_nl));
  assign ACCUM_INNER_LOOP_1_acc_140_nl = nl_ACCUM_INNER_LOOP_1_acc_140_nl[15:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_328_0}))
      * $signed((w5_rsci_idat[1749:1745]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_330_0}))
      * $signed((w5_rsci_idat[1734:1730]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_320_0}))
      * $signed((w5_rsci_idat[1769:1765]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_322_0}))
      * $signed((w5_rsci_idat[1754:1750]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_344_0}))
      * $signed((w5_rsci_idat[1709:1705]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_346_0}))
      * $signed((w5_rsci_idat[1694:1690]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_336_0}))
      * $signed((w5_rsci_idat[1729:1725]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_338_0}))
      * $signed((w5_rsci_idat[1714:1710]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_340_0}))
      * $signed((w5_rsci_idat[1719:1715]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_342_0}))
      * $signed((w5_rsci_idat[1704:1700]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_352_0}))
      * $signed((w5_rsci_idat[1689:1685]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_354_0}))
      * $signed((w5_rsci_idat[1674:1670]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_356_0}))
      * $signed((w5_rsci_idat[1679:1675]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_358_0}))
      * $signed((w5_rsci_idat[1664:1660]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_360_0}))
      * $signed((w5_rsci_idat[1669:1665]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_362_0}))
      * $signed((w5_rsci_idat[1654:1650]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_364_0}))
      * $signed((w5_rsci_idat[1659:1655]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_366_0}))
      * $signed((w5_rsci_idat[1644:1640]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_376_0}))
      * $signed((w5_rsci_idat[1629:1625]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_378_0}))
      * $signed((w5_rsci_idat[1614:1610]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_380_0}))
      * $signed((w5_rsci_idat[1619:1615]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_382_0}))
      * $signed((w5_rsci_idat[1604:1600]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_368_0}))
      * $signed((w5_rsci_idat[1649:1645]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_370_0}))
      * $signed((w5_rsci_idat[1634:1630]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_372_0}))
      * $signed((w5_rsci_idat[1639:1635]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_374_0}))
      * $signed((w5_rsci_idat[1624:1620]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_324_0}))
      * $signed((w5_rsci_idat[1759:1755]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_326_0}))
      * $signed((w5_rsci_idat[1744:1740]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_332_0}))
      * $signed((w5_rsci_idat[1739:1735]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_334_0}))
      * $signed((w5_rsci_idat[1724:1720]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_348_0}))
      * $signed((w5_rsci_idat[1699:1695]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_9
      , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_8_1 , nnet_relu_layer2_t_layer4_t_relu_config4_for_if_conc_350_0}))
      * $signed((w5_rsci_idat[1684:1680]));
  assign ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl = nl_ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl[14:0];
  assign nl_layer5_out_rsci_idat_47_32  = ACCUM_INNER_LOOP_1_acc_139_nl + ACCUM_INNER_LOOP_1_acc_140_nl
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_94_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_91_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_98_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_95_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_86_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_83_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_90_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_87_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_88_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_85_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_82_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_79_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_80_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_77_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_78_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_75_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_76_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_73_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_70_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_67_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_68_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_65_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_74_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_71_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_72_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_69_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_96_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_93_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_92_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_89_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_84_ACCUM_INNER_LOOP_1_mul_nl))
      + conv_s2s_11_16(readslicef_15_11_4(ACCUM_OUTER_LOOP_1_3_ACCUM_INNER_LOOP_1_81_ACCUM_INNER_LOOP_1_mul_nl));

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [10:0] readslicef_15_11_4;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_15_11_4 = tmp[10:0];
  end
  endfunction


  function automatic [0:0] readslicef_17_1_16;
    input [16:0] vector;
    reg [16:0] tmp;
  begin
    tmp = vector >> 16;
    readslicef_17_1_16 = tmp[0:0];
  end
  endfunction


  function automatic [15:0] readslicef_20_16_4;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_20_16_4 = tmp[15:0];
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_5_10 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_10 = {{5{vector[4]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_11_16 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_16 = {{5{vector[10]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_12_16 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_16 = {{4{vector[11]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    myproject
// ------------------------------------------------------------------


module myproject (
  clk, rst, input_1_rsc_dat, layer5_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [223:0] input_1_rsc_dat;
  output [47:0] layer5_out_rsc_dat;
  input [8959:0] w2_rsc_dat;
  input [639:0] b2_rsc_dat;
  input [1919:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  converterBlock_myproject_core myproject_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .w2_rsc_dat(w2_rsc_dat),
      .b2_rsc_dat(b2_rsc_dat),
      .w5_rsc_dat(w5_rsc_dat),
      .b5_rsc_dat(b5_rsc_dat)
    );
endmodule



