
//------> ./myproject_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module converterBlock_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./myproject_ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module converterBlock_ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./myproject.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
// 
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Mon Feb 13 21:34:31 2023
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core
// ------------------------------------------------------------------


module converterBlock_myproject_core (
  clk, rst, input_1_rsc_dat, layer7_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [95:0] input_1_rsc_dat;
  output [1:0] layer7_out_rsc_dat;
  input [4639:0] w2_rsc_dat;
  input [289:0] b2_rsc_dat;
  input [869:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;


  // Interconnect Declarations
  wire [95:0] input_1_rsci_idat;
  reg [1:0] layer7_out_rsci_idat;
  wire [4639:0] w2_rsci_idat;
  wire [289:0] b2_rsci_idat;
  wire [869:0] w5_rsci_idat;
  wire [14:0] b5_rsci_idat;
  wire [8:0] Accum2_acc_121_psp_sva_1;
  wire [9:0] nl_Accum2_acc_121_psp_sva_1;
  wire [8:0] Accum2_acc_120_psp_sva_1;
  wire [9:0] nl_Accum2_acc_120_psp_sva_1;
  wire [8:0] Accum2_acc_119_psp_sva_1;
  wire [9:0] nl_Accum2_acc_119_psp_sva_1;
  wire [8:0] Accum2_acc_118_psp_sva_1;
  wire [9:0] nl_Accum2_acc_118_psp_sva_1;
  wire [8:0] Accum2_acc_117_psp_sva_1;
  wire [9:0] nl_Accum2_acc_117_psp_sva_1;
  wire [8:0] Accum2_acc_116_psp_sva_1;
  wire [9:0] nl_Accum2_acc_116_psp_sva_1;
  wire [8:0] Accum2_acc_115_psp_sva_1;
  wire [9:0] nl_Accum2_acc_115_psp_sva_1;
  wire [8:0] Accum2_acc_114_psp_sva_1;
  wire [9:0] nl_Accum2_acc_114_psp_sva_1;
  wire [8:0] Accum2_acc_113_psp_sva_1;
  wire [9:0] nl_Accum2_acc_113_psp_sva_1;
  wire [8:0] Accum2_acc_112_psp_sva_1;
  wire [9:0] nl_Accum2_acc_112_psp_sva_1;
  wire [8:0] Accum2_acc_111_psp_sva_1;
  wire [9:0] nl_Accum2_acc_111_psp_sva_1;
  wire [8:0] Accum2_acc_110_psp_sva_1;
  wire [9:0] nl_Accum2_acc_110_psp_sva_1;
  wire [8:0] Accum2_acc_109_psp_sva_1;
  wire [9:0] nl_Accum2_acc_109_psp_sva_1;
  wire [8:0] Accum2_acc_108_psp_sva_1;
  wire [9:0] nl_Accum2_acc_108_psp_sva_1;
  wire [8:0] Accum2_acc_107_psp_sva_1;
  wire [9:0] nl_Accum2_acc_107_psp_sva_1;
  wire [8:0] Accum2_acc_106_psp_sva_1;
  wire [9:0] nl_Accum2_acc_106_psp_sva_1;
  wire [8:0] Accum2_acc_105_psp_sva_1;
  wire [9:0] nl_Accum2_acc_105_psp_sva_1;
  wire [8:0] Accum2_acc_104_psp_sva_1;
  wire [9:0] nl_Accum2_acc_104_psp_sva_1;
  wire [8:0] Accum2_acc_103_psp_sva_1;
  wire [9:0] nl_Accum2_acc_103_psp_sva_1;
  wire [8:0] Accum2_acc_102_psp_sva_1;
  wire [9:0] nl_Accum2_acc_102_psp_sva_1;
  wire [8:0] Accum2_acc_101_psp_sva_1;
  wire [9:0] nl_Accum2_acc_101_psp_sva_1;
  wire [8:0] Accum2_acc_100_psp_sva_1;
  wire [9:0] nl_Accum2_acc_100_psp_sva_1;
  wire [8:0] Accum2_acc_99_psp_sva_1;
  wire [9:0] nl_Accum2_acc_99_psp_sva_1;
  wire [8:0] Accum2_acc_98_psp_sva_1;
  wire [9:0] nl_Accum2_acc_98_psp_sva_1;
  wire [8:0] Accum2_acc_97_psp_sva_1;
  wire [9:0] nl_Accum2_acc_97_psp_sva_1;
  wire [8:0] Accum2_acc_96_psp_sva_1;
  wire [9:0] nl_Accum2_acc_96_psp_sva_1;
  wire [8:0] Accum2_acc_95_psp_sva_1;
  wire [9:0] nl_Accum2_acc_95_psp_sva_1;
  wire [8:0] Accum2_acc_94_psp_sva_1;
  wire [9:0] nl_Accum2_acc_94_psp_sva_1;
  wire [8:0] Accum2_acc_93_psp_sva_1;
  wire [9:0] nl_Accum2_acc_93_psp_sva_1;
  wire [8:0] Accum2_acc_92_psp_sva_1;
  wire [9:0] nl_Accum2_acc_92_psp_sva_1;
  wire [8:0] Accum2_acc_91_psp_sva_1;
  wire [9:0] nl_Accum2_acc_91_psp_sva_1;
  wire [8:0] Accum2_acc_90_psp_sva_1;
  wire [9:0] nl_Accum2_acc_90_psp_sva_1;
  wire [8:0] Accum2_acc_89_psp_sva_1;
  wire [9:0] nl_Accum2_acc_89_psp_sva_1;
  wire [8:0] Accum2_acc_88_psp_sva_1;
  wire [9:0] nl_Accum2_acc_88_psp_sva_1;
  wire [8:0] Accum2_acc_87_psp_sva_1;
  wire [9:0] nl_Accum2_acc_87_psp_sva_1;
  wire [8:0] Accum2_acc_86_psp_sva_1;
  wire [9:0] nl_Accum2_acc_86_psp_sva_1;
  wire [8:0] Accum2_acc_85_psp_sva_1;
  wire [9:0] nl_Accum2_acc_85_psp_sva_1;
  wire [8:0] Accum2_acc_84_psp_sva_1;
  wire [9:0] nl_Accum2_acc_84_psp_sva_1;
  wire [8:0] Accum2_acc_83_psp_sva_1;
  wire [9:0] nl_Accum2_acc_83_psp_sva_1;
  wire [8:0] Accum2_acc_82_psp_sva_1;
  wire [9:0] nl_Accum2_acc_82_psp_sva_1;
  wire [8:0] Accum2_acc_81_psp_sva_1;
  wire [9:0] nl_Accum2_acc_81_psp_sva_1;
  wire [8:0] Accum2_acc_80_psp_sva_1;
  wire [9:0] nl_Accum2_acc_80_psp_sva_1;
  wire [8:0] Accum2_acc_79_psp_sva_1;
  wire [9:0] nl_Accum2_acc_79_psp_sva_1;
  wire [8:0] Accum2_acc_78_psp_sva_1;
  wire [9:0] nl_Accum2_acc_78_psp_sva_1;
  wire [8:0] Accum2_acc_77_psp_sva_1;
  wire [9:0] nl_Accum2_acc_77_psp_sva_1;
  wire [8:0] Accum2_acc_76_psp_sva_1;
  wire [9:0] nl_Accum2_acc_76_psp_sva_1;
  wire [8:0] Accum2_acc_75_psp_sva_1;
  wire [9:0] nl_Accum2_acc_75_psp_sva_1;
  wire [8:0] Accum2_acc_74_psp_sva_1;
  wire [9:0] nl_Accum2_acc_74_psp_sva_1;
  wire [8:0] Accum2_acc_73_psp_sva_1;
  wire [9:0] nl_Accum2_acc_73_psp_sva_1;
  wire [8:0] Accum2_acc_72_psp_sva_1;
  wire [9:0] nl_Accum2_acc_72_psp_sva_1;
  wire [8:0] Accum2_acc_71_psp_sva_1;
  wire [9:0] nl_Accum2_acc_71_psp_sva_1;
  wire [8:0] Accum2_acc_70_psp_sva_1;
  wire [9:0] nl_Accum2_acc_70_psp_sva_1;
  wire [8:0] Accum2_acc_69_psp_sva_1;
  wire [9:0] nl_Accum2_acc_69_psp_sva_1;
  wire [8:0] Accum2_acc_68_psp_sva_1;
  wire [9:0] nl_Accum2_acc_68_psp_sva_1;
  wire [8:0] Accum2_acc_67_psp_sva_1;
  wire [9:0] nl_Accum2_acc_67_psp_sva_1;
  wire [8:0] Accum2_acc_66_psp_sva_1;
  wire [9:0] nl_Accum2_acc_66_psp_sva_1;
  wire [8:0] Accum2_acc_65_psp_sva_1;
  wire [9:0] nl_Accum2_acc_65_psp_sva_1;
  wire [8:0] layer3_out_0_9_1_sva_1;
  wire [9:0] nl_layer3_out_0_9_1_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire layer4_out_0_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_8_6;
  wire layer4_out_conc_4_9;
  wire [2:0] layer4_out_conc_4_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_8_6;
  wire [9:0] Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_itm_12_3_1;
  wire [9:0] Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_itm_12_3_1;
  wire [9:0] Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_itm_12_3_1;
  wire [8:0] Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1;
  wire [8:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1;
  wire [8:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;

  wire[1:0] argmax_else_mux_nl;
  wire argmax_else_if_argmax_else_if_argmax_else_if_nor_nl;
  wire[10:0] argmax_else_aif_acc_nl;
  wire[11:0] nl_argmax_else_aif_acc_nl;
  wire[10:0] argmax_else_acc_nl;
  wire[11:0] nl_argmax_else_acc_nl;
  wire argmax_if_argmax_if_argmax_if_nor_nl;
  wire[10:0] argmax_aif_acc_nl;
  wire[11:0] nl_argmax_aif_acc_nl;
  wire[10:0] argmax_acc_nl;
  wire[11:0] nl_argmax_acc_nl;
  wire[8:0] Accum2_acc_1782_nl;
  wire[9:0] nl_Accum2_acc_1782_nl;
  wire[8:0] Accum2_acc_1780_nl;
  wire[9:0] nl_Accum2_acc_1780_nl;
  wire[8:0] Accum2_acc_1776_nl;
  wire[9:0] nl_Accum2_acc_1776_nl;
  wire[8:0] Accum2_acc_1768_nl;
  wire[9:0] nl_Accum2_acc_1768_nl;
  wire[8:0] Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1775_nl;
  wire[9:0] nl_Accum2_acc_1775_nl;
  wire[8:0] Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1779_nl;
  wire[10:0] nl_Accum2_acc_1779_nl;
  wire[8:0] Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1781_nl;
  wire[11:0] nl_Accum2_acc_1781_nl;
  wire[8:0] Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_nl;
  wire[11:0] nl_Accum2_acc_nl;
  wire[8:0] Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_921_nl;
  wire[9:0] nl_Accum2_acc_921_nl;
  wire[8:0] Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_926_nl;
  wire[11:0] nl_Accum2_acc_926_nl;
  wire[8:0] Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_942_nl;
  wire[11:0] nl_Accum2_acc_942_nl;
  wire[8:0] Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_928_nl;
  wire[9:0] nl_Accum2_acc_928_nl;
  wire[8:0] Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_941_nl;
  wire[11:0] nl_Accum2_acc_941_nl;
  wire[8:0] Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_957_nl;
  wire[11:0] nl_Accum2_acc_957_nl;
  wire[8:0] Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_943_nl;
  wire[9:0] nl_Accum2_acc_943_nl;
  wire[8:0] Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_956_nl;
  wire[11:0] nl_Accum2_acc_956_nl;
  wire[8:0] Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_972_nl;
  wire[11:0] nl_Accum2_acc_972_nl;
  wire[8:0] Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_958_nl;
  wire[9:0] nl_Accum2_acc_958_nl;
  wire[8:0] Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_971_nl;
  wire[11:0] nl_Accum2_acc_971_nl;
  wire[8:0] Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_987_nl;
  wire[11:0] nl_Accum2_acc_987_nl;
  wire[8:0] Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_973_nl;
  wire[9:0] nl_Accum2_acc_973_nl;
  wire[8:0] Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_986_nl;
  wire[11:0] nl_Accum2_acc_986_nl;
  wire[8:0] Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1002_nl;
  wire[11:0] nl_Accum2_acc_1002_nl;
  wire[8:0] Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_988_nl;
  wire[9:0] nl_Accum2_acc_988_nl;
  wire[8:0] Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1001_nl;
  wire[11:0] nl_Accum2_acc_1001_nl;
  wire[8:0] Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1017_nl;
  wire[11:0] nl_Accum2_acc_1017_nl;
  wire[8:0] Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1003_nl;
  wire[9:0] nl_Accum2_acc_1003_nl;
  wire[8:0] Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1016_nl;
  wire[11:0] nl_Accum2_acc_1016_nl;
  wire[8:0] Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1032_nl;
  wire[11:0] nl_Accum2_acc_1032_nl;
  wire[8:0] Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1018_nl;
  wire[9:0] nl_Accum2_acc_1018_nl;
  wire[8:0] Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1031_nl;
  wire[11:0] nl_Accum2_acc_1031_nl;
  wire[8:0] Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1047_nl;
  wire[11:0] nl_Accum2_acc_1047_nl;
  wire[8:0] Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1033_nl;
  wire[9:0] nl_Accum2_acc_1033_nl;
  wire[8:0] Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1046_nl;
  wire[11:0] nl_Accum2_acc_1046_nl;
  wire[8:0] Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1062_nl;
  wire[11:0] nl_Accum2_acc_1062_nl;
  wire[8:0] Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1048_nl;
  wire[9:0] nl_Accum2_acc_1048_nl;
  wire[8:0] Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1061_nl;
  wire[11:0] nl_Accum2_acc_1061_nl;
  wire[8:0] Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1077_nl;
  wire[11:0] nl_Accum2_acc_1077_nl;
  wire[8:0] Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1063_nl;
  wire[9:0] nl_Accum2_acc_1063_nl;
  wire[8:0] Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1076_nl;
  wire[11:0] nl_Accum2_acc_1076_nl;
  wire[8:0] Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1092_nl;
  wire[11:0] nl_Accum2_acc_1092_nl;
  wire[8:0] Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1078_nl;
  wire[9:0] nl_Accum2_acc_1078_nl;
  wire[8:0] Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1091_nl;
  wire[11:0] nl_Accum2_acc_1091_nl;
  wire[8:0] Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1107_nl;
  wire[11:0] nl_Accum2_acc_1107_nl;
  wire[8:0] Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1093_nl;
  wire[9:0] nl_Accum2_acc_1093_nl;
  wire[8:0] Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1106_nl;
  wire[11:0] nl_Accum2_acc_1106_nl;
  wire[8:0] Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1122_nl;
  wire[11:0] nl_Accum2_acc_1122_nl;
  wire[8:0] Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1108_nl;
  wire[9:0] nl_Accum2_acc_1108_nl;
  wire[8:0] Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1121_nl;
  wire[11:0] nl_Accum2_acc_1121_nl;
  wire[8:0] Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1137_nl;
  wire[11:0] nl_Accum2_acc_1137_nl;
  wire[8:0] Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1123_nl;
  wire[9:0] nl_Accum2_acc_1123_nl;
  wire[8:0] Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1136_nl;
  wire[11:0] nl_Accum2_acc_1136_nl;
  wire[8:0] Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1152_nl;
  wire[11:0] nl_Accum2_acc_1152_nl;
  wire[8:0] Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1138_nl;
  wire[9:0] nl_Accum2_acc_1138_nl;
  wire[8:0] Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1151_nl;
  wire[11:0] nl_Accum2_acc_1151_nl;
  wire[8:0] Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1167_nl;
  wire[11:0] nl_Accum2_acc_1167_nl;
  wire[8:0] Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1153_nl;
  wire[9:0] nl_Accum2_acc_1153_nl;
  wire[8:0] Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1166_nl;
  wire[11:0] nl_Accum2_acc_1166_nl;
  wire[8:0] Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1182_nl;
  wire[11:0] nl_Accum2_acc_1182_nl;
  wire[8:0] Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1168_nl;
  wire[9:0] nl_Accum2_acc_1168_nl;
  wire[8:0] Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1181_nl;
  wire[11:0] nl_Accum2_acc_1181_nl;
  wire[8:0] Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1197_nl;
  wire[11:0] nl_Accum2_acc_1197_nl;
  wire[8:0] Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1183_nl;
  wire[9:0] nl_Accum2_acc_1183_nl;
  wire[8:0] Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1196_nl;
  wire[11:0] nl_Accum2_acc_1196_nl;
  wire[8:0] Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1212_nl;
  wire[11:0] nl_Accum2_acc_1212_nl;
  wire[8:0] Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1198_nl;
  wire[9:0] nl_Accum2_acc_1198_nl;
  wire[8:0] Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1211_nl;
  wire[11:0] nl_Accum2_acc_1211_nl;
  wire[8:0] Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1227_nl;
  wire[11:0] nl_Accum2_acc_1227_nl;
  wire[8:0] Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1213_nl;
  wire[9:0] nl_Accum2_acc_1213_nl;
  wire[8:0] Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1226_nl;
  wire[11:0] nl_Accum2_acc_1226_nl;
  wire[8:0] Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1242_nl;
  wire[11:0] nl_Accum2_acc_1242_nl;
  wire[8:0] Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1228_nl;
  wire[9:0] nl_Accum2_acc_1228_nl;
  wire[8:0] Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1241_nl;
  wire[11:0] nl_Accum2_acc_1241_nl;
  wire[8:0] Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1257_nl;
  wire[11:0] nl_Accum2_acc_1257_nl;
  wire[8:0] Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1243_nl;
  wire[9:0] nl_Accum2_acc_1243_nl;
  wire[8:0] Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1256_nl;
  wire[11:0] nl_Accum2_acc_1256_nl;
  wire[8:0] Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1272_nl;
  wire[11:0] nl_Accum2_acc_1272_nl;
  wire[8:0] Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1258_nl;
  wire[9:0] nl_Accum2_acc_1258_nl;
  wire[8:0] Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1271_nl;
  wire[11:0] nl_Accum2_acc_1271_nl;
  wire[8:0] Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1287_nl;
  wire[11:0] nl_Accum2_acc_1287_nl;
  wire[8:0] Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1273_nl;
  wire[9:0] nl_Accum2_acc_1273_nl;
  wire[8:0] Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1286_nl;
  wire[11:0] nl_Accum2_acc_1286_nl;
  wire[8:0] Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1302_nl;
  wire[11:0] nl_Accum2_acc_1302_nl;
  wire[8:0] Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1288_nl;
  wire[9:0] nl_Accum2_acc_1288_nl;
  wire[8:0] Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1301_nl;
  wire[11:0] nl_Accum2_acc_1301_nl;
  wire[8:0] Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1317_nl;
  wire[11:0] nl_Accum2_acc_1317_nl;
  wire[8:0] Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1303_nl;
  wire[9:0] nl_Accum2_acc_1303_nl;
  wire[8:0] Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1316_nl;
  wire[11:0] nl_Accum2_acc_1316_nl;
  wire[8:0] Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1332_nl;
  wire[11:0] nl_Accum2_acc_1332_nl;
  wire[8:0] Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1318_nl;
  wire[9:0] nl_Accum2_acc_1318_nl;
  wire[8:0] Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1331_nl;
  wire[11:0] nl_Accum2_acc_1331_nl;
  wire[8:0] Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1347_nl;
  wire[11:0] nl_Accum2_acc_1347_nl;
  wire[8:0] Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1333_nl;
  wire[9:0] nl_Accum2_acc_1333_nl;
  wire[8:0] Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1346_nl;
  wire[11:0] nl_Accum2_acc_1346_nl;
  wire[8:0] Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1362_nl;
  wire[11:0] nl_Accum2_acc_1362_nl;
  wire[8:0] Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1348_nl;
  wire[9:0] nl_Accum2_acc_1348_nl;
  wire[8:0] Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1361_nl;
  wire[11:0] nl_Accum2_acc_1361_nl;
  wire[8:0] Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1377_nl;
  wire[11:0] nl_Accum2_acc_1377_nl;
  wire[8:0] Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1363_nl;
  wire[9:0] nl_Accum2_acc_1363_nl;
  wire[8:0] Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1376_nl;
  wire[11:0] nl_Accum2_acc_1376_nl;
  wire[8:0] Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1392_nl;
  wire[11:0] nl_Accum2_acc_1392_nl;
  wire[8:0] Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1378_nl;
  wire[9:0] nl_Accum2_acc_1378_nl;
  wire[8:0] Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1391_nl;
  wire[11:0] nl_Accum2_acc_1391_nl;
  wire[8:0] Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1407_nl;
  wire[11:0] nl_Accum2_acc_1407_nl;
  wire[8:0] Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1393_nl;
  wire[9:0] nl_Accum2_acc_1393_nl;
  wire[8:0] Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1406_nl;
  wire[11:0] nl_Accum2_acc_1406_nl;
  wire[8:0] Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1422_nl;
  wire[11:0] nl_Accum2_acc_1422_nl;
  wire[8:0] Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1408_nl;
  wire[9:0] nl_Accum2_acc_1408_nl;
  wire[8:0] Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1421_nl;
  wire[11:0] nl_Accum2_acc_1421_nl;
  wire[8:0] Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1437_nl;
  wire[11:0] nl_Accum2_acc_1437_nl;
  wire[8:0] Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1423_nl;
  wire[9:0] nl_Accum2_acc_1423_nl;
  wire[8:0] Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1436_nl;
  wire[11:0] nl_Accum2_acc_1436_nl;
  wire[8:0] Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1452_nl;
  wire[11:0] nl_Accum2_acc_1452_nl;
  wire[8:0] Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1438_nl;
  wire[9:0] nl_Accum2_acc_1438_nl;
  wire[8:0] Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1451_nl;
  wire[11:0] nl_Accum2_acc_1451_nl;
  wire[8:0] Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1467_nl;
  wire[11:0] nl_Accum2_acc_1467_nl;
  wire[8:0] Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1453_nl;
  wire[9:0] nl_Accum2_acc_1453_nl;
  wire[8:0] Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1466_nl;
  wire[11:0] nl_Accum2_acc_1466_nl;
  wire[8:0] Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1482_nl;
  wire[11:0] nl_Accum2_acc_1482_nl;
  wire[8:0] Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1468_nl;
  wire[9:0] nl_Accum2_acc_1468_nl;
  wire[8:0] Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1481_nl;
  wire[11:0] nl_Accum2_acc_1481_nl;
  wire[8:0] Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1497_nl;
  wire[11:0] nl_Accum2_acc_1497_nl;
  wire[8:0] Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1483_nl;
  wire[9:0] nl_Accum2_acc_1483_nl;
  wire[8:0] Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1496_nl;
  wire[11:0] nl_Accum2_acc_1496_nl;
  wire[8:0] Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1512_nl;
  wire[11:0] nl_Accum2_acc_1512_nl;
  wire[8:0] Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1498_nl;
  wire[9:0] nl_Accum2_acc_1498_nl;
  wire[8:0] Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1511_nl;
  wire[11:0] nl_Accum2_acc_1511_nl;
  wire[8:0] Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1527_nl;
  wire[11:0] nl_Accum2_acc_1527_nl;
  wire[8:0] Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1513_nl;
  wire[9:0] nl_Accum2_acc_1513_nl;
  wire[8:0] Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1526_nl;
  wire[11:0] nl_Accum2_acc_1526_nl;
  wire[8:0] Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1542_nl;
  wire[11:0] nl_Accum2_acc_1542_nl;
  wire[8:0] Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1528_nl;
  wire[9:0] nl_Accum2_acc_1528_nl;
  wire[8:0] Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1541_nl;
  wire[11:0] nl_Accum2_acc_1541_nl;
  wire[8:0] Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1557_nl;
  wire[11:0] nl_Accum2_acc_1557_nl;
  wire[8:0] Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1543_nl;
  wire[9:0] nl_Accum2_acc_1543_nl;
  wire[8:0] Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1556_nl;
  wire[11:0] nl_Accum2_acc_1556_nl;
  wire[8:0] Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1572_nl;
  wire[11:0] nl_Accum2_acc_1572_nl;
  wire[8:0] Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1558_nl;
  wire[9:0] nl_Accum2_acc_1558_nl;
  wire[8:0] Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1571_nl;
  wire[11:0] nl_Accum2_acc_1571_nl;
  wire[8:0] Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1587_nl;
  wire[11:0] nl_Accum2_acc_1587_nl;
  wire[8:0] Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1573_nl;
  wire[9:0] nl_Accum2_acc_1573_nl;
  wire[8:0] Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1586_nl;
  wire[11:0] nl_Accum2_acc_1586_nl;
  wire[8:0] Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1602_nl;
  wire[11:0] nl_Accum2_acc_1602_nl;
  wire[8:0] Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1588_nl;
  wire[9:0] nl_Accum2_acc_1588_nl;
  wire[8:0] Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1601_nl;
  wire[11:0] nl_Accum2_acc_1601_nl;
  wire[8:0] Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1617_nl;
  wire[11:0] nl_Accum2_acc_1617_nl;
  wire[8:0] Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1603_nl;
  wire[9:0] nl_Accum2_acc_1603_nl;
  wire[8:0] Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1616_nl;
  wire[11:0] nl_Accum2_acc_1616_nl;
  wire[8:0] Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1632_nl;
  wire[11:0] nl_Accum2_acc_1632_nl;
  wire[8:0] Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1618_nl;
  wire[9:0] nl_Accum2_acc_1618_nl;
  wire[8:0] Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1631_nl;
  wire[11:0] nl_Accum2_acc_1631_nl;
  wire[8:0] Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1647_nl;
  wire[11:0] nl_Accum2_acc_1647_nl;
  wire[8:0] Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1633_nl;
  wire[9:0] nl_Accum2_acc_1633_nl;
  wire[8:0] Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1646_nl;
  wire[11:0] nl_Accum2_acc_1646_nl;
  wire[8:0] Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1662_nl;
  wire[11:0] nl_Accum2_acc_1662_nl;
  wire[8:0] Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1648_nl;
  wire[9:0] nl_Accum2_acc_1648_nl;
  wire[8:0] Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1661_nl;
  wire[11:0] nl_Accum2_acc_1661_nl;
  wire[8:0] Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1677_nl;
  wire[11:0] nl_Accum2_acc_1677_nl;
  wire[8:0] Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1663_nl;
  wire[9:0] nl_Accum2_acc_1663_nl;
  wire[8:0] Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1676_nl;
  wire[11:0] nl_Accum2_acc_1676_nl;
  wire[8:0] Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1692_nl;
  wire[11:0] nl_Accum2_acc_1692_nl;
  wire[8:0] Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1678_nl;
  wire[9:0] nl_Accum2_acc_1678_nl;
  wire[8:0] Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1691_nl;
  wire[11:0] nl_Accum2_acc_1691_nl;
  wire[8:0] Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1707_nl;
  wire[11:0] nl_Accum2_acc_1707_nl;
  wire[8:0] Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1693_nl;
  wire[9:0] nl_Accum2_acc_1693_nl;
  wire[8:0] Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1706_nl;
  wire[11:0] nl_Accum2_acc_1706_nl;
  wire[8:0] Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1722_nl;
  wire[11:0] nl_Accum2_acc_1722_nl;
  wire[8:0] Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1708_nl;
  wire[9:0] nl_Accum2_acc_1708_nl;
  wire[8:0] Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1721_nl;
  wire[11:0] nl_Accum2_acc_1721_nl;
  wire[8:0] Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1737_nl;
  wire[11:0] nl_Accum2_acc_1737_nl;
  wire[8:0] Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1723_nl;
  wire[9:0] nl_Accum2_acc_1723_nl;
  wire[8:0] Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1736_nl;
  wire[11:0] nl_Accum2_acc_1736_nl;
  wire[8:0] Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1752_nl;
  wire[11:0] nl_Accum2_acc_1752_nl;
  wire[8:0] Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1738_nl;
  wire[9:0] nl_Accum2_acc_1738_nl;
  wire[8:0] Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1751_nl;
  wire[11:0] nl_Accum2_acc_1751_nl;
  wire[8:0] Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1767_nl;
  wire[11:0] nl_Accum2_acc_1767_nl;
  wire[8:0] Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1753_nl;
  wire[9:0] nl_Accum2_acc_1753_nl;
  wire[8:0] Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Accum2_acc_1766_nl;
  wire[11:0] nl_Accum2_acc_1766_nl;
  wire[8:0] Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[8:0] Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[12:0] Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_nl;
  wire[17:0] nl_Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_nl;
  wire[12:0] Accum2_1_acc_114_nl;
  wire[17:0] nl_Accum2_1_acc_114_nl;
  wire[14:0] Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_174_nl;
  wire[6:0] nl_Accum2_1_acc_174_nl;
  wire[14:0] Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[12:0] Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_nl;
  wire[17:0] nl_Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_nl;
  wire[12:0] Accum2_1_acc_171_nl;
  wire[17:0] nl_Accum2_1_acc_171_nl;
  wire[14:0] Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_175_nl;
  wire[6:0] nl_Accum2_1_acc_175_nl;
  wire[14:0] Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[12:0] Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_nl;
  wire[17:0] nl_Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_nl;
  wire[12:0] Accum2_1_acc_nl;
  wire[17:0] nl_Accum2_1_acc_nl;
  wire[14:0] Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_173_nl;
  wire[6:0] nl_Accum2_1_acc_173_nl;
  wire[14:0] Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[10:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[11:0] nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;

  // Interconnect Declarations for Component Instantiations 
  converterBlock_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd96)) input_1_rsci (
      .dat(input_1_rsc_dat),
      .idat(input_1_rsci_idat)
    );
  converterBlock_ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd2)) layer7_out_rsci (
      .idat(layer7_out_rsci_idat),
      .dat(layer7_out_rsc_dat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd4640)) w2_rsci (
      .dat(w2_rsc_dat),
      .idat(w2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd290)) b2_rsci (
      .dat(b2_rsc_dat),
      .idat(b2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd870)) w5_rsci (
      .dat(w5_rsc_dat),
      .idat(w5_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd15)) b5_rsci (
      .dat(b5_rsc_dat),
      .idat(b5_rsci_idat)
    );
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1 = (layer3_out_0_9_1_sva_1[7:4]!=4'b0000);
  assign nl_Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4354:4350]));
  assign Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1768_nl = Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[4:0]);
  assign Accum2_acc_1768_nl = nl_Accum2_acc_1768_nl[8:0];
  assign nl_Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[4:0]));
  assign Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1776_nl = Accum2_acc_1768_nl + Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1776_nl = nl_Accum2_acc_1776_nl[8:0];
  assign nl_Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[294:290]));
  assign Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[584:580]));
  assign Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1775_nl = Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1775_nl = nl_Accum2_acc_1775_nl[8:0];
  assign nl_Accum2_acc_1780_nl = Accum2_acc_1776_nl + Accum2_acc_1775_nl;
  assign Accum2_acc_1780_nl = nl_Accum2_acc_1780_nl[8:0];
  assign nl_Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[874:870]));
  assign Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1164:1160]));
  assign Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1454:1450]));
  assign Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1744:1740]));
  assign Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1779_nl = Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1779_nl = nl_Accum2_acc_1779_nl[8:0];
  assign nl_Accum2_acc_1782_nl = Accum2_acc_1780_nl + Accum2_acc_1779_nl;
  assign Accum2_acc_1782_nl = nl_Accum2_acc_1782_nl[8:0];
  assign nl_Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3194:3190]));
  assign Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3484:3480]));
  assign Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2034:2030]));
  assign Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2324:2320]));
  assign Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2614:2610]));
  assign Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2904:2900]));
  assign Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3774:3770]));
  assign Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4064:4060]));
  assign Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1781_nl = Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1781_nl = nl_Accum2_acc_1781_nl[8:0];
  assign nl_layer3_out_0_9_1_sva_1 = Accum2_acc_1782_nl + Accum2_acc_1781_nl;
  assign layer3_out_0_9_1_sva_1 = nl_layer3_out_0_9_1_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 = (Accum2_acc_65_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[879:875]));
  assign Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1169:1165]));
  assign Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4359:4355]));
  assign Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_921_nl = Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[9:5]);
  assign Accum2_acc_921_nl = nl_Accum2_acc_921_nl[8:0];
  assign nl_Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[9:5]));
  assign Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[299:295]));
  assign Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[589:585]));
  assign Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1459:1455]));
  assign Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1749:1745]));
  assign Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_nl = Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_921_nl
      + Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_nl = nl_Accum2_acc_nl[8:0];
  assign nl_Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3199:3195]));
  assign Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3489:3485]));
  assign Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2039:2035]));
  assign Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2329:2325]));
  assign Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2619:2615]));
  assign Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2909:2905]));
  assign Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3779:3775]));
  assign Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4069:4065]));
  assign Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_926_nl = Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_926_nl = nl_Accum2_acc_926_nl[8:0];
  assign nl_Accum2_acc_65_psp_sva_1 = Accum2_acc_nl + Accum2_acc_926_nl;
  assign Accum2_acc_65_psp_sva_1 = nl_Accum2_acc_65_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 = (Accum2_acc_66_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[884:880]));
  assign Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1174:1170]));
  assign Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4364:4360]));
  assign Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_928_nl = Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[14:10]);
  assign Accum2_acc_928_nl = nl_Accum2_acc_928_nl[8:0];
  assign nl_Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[14:10]));
  assign Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[304:300]));
  assign Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[594:590]));
  assign Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1464:1460]));
  assign Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1754:1750]));
  assign Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_942_nl = Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_928_nl
      + Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_942_nl = nl_Accum2_acc_942_nl[8:0];
  assign nl_Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3204:3200]));
  assign Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3494:3490]));
  assign Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2044:2040]));
  assign Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2334:2330]));
  assign Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2624:2620]));
  assign Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2914:2910]));
  assign Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3784:3780]));
  assign Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4074:4070]));
  assign Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_941_nl = Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_941_nl = nl_Accum2_acc_941_nl[8:0];
  assign nl_Accum2_acc_66_psp_sva_1 = Accum2_acc_942_nl + Accum2_acc_941_nl;
  assign Accum2_acc_66_psp_sva_1 = nl_Accum2_acc_66_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 = (Accum2_acc_67_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[889:885]));
  assign Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1179:1175]));
  assign Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4369:4365]));
  assign Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_943_nl = Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[19:15]);
  assign Accum2_acc_943_nl = nl_Accum2_acc_943_nl[8:0];
  assign nl_Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[19:15]));
  assign Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[309:305]));
  assign Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[599:595]));
  assign Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1469:1465]));
  assign Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1759:1755]));
  assign Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_957_nl = Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_943_nl
      + Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_957_nl = nl_Accum2_acc_957_nl[8:0];
  assign nl_Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3209:3205]));
  assign Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3499:3495]));
  assign Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2049:2045]));
  assign Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2339:2335]));
  assign Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2629:2625]));
  assign Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2919:2915]));
  assign Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3789:3785]));
  assign Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4079:4075]));
  assign Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_956_nl = Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_956_nl = nl_Accum2_acc_956_nl[8:0];
  assign nl_Accum2_acc_67_psp_sva_1 = Accum2_acc_957_nl + Accum2_acc_956_nl;
  assign Accum2_acc_67_psp_sva_1 = nl_Accum2_acc_67_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 = (Accum2_acc_68_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[894:890]));
  assign Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1184:1180]));
  assign Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4374:4370]));
  assign Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_958_nl = Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[24:20]);
  assign Accum2_acc_958_nl = nl_Accum2_acc_958_nl[8:0];
  assign nl_Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[24:20]));
  assign Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[314:310]));
  assign Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[604:600]));
  assign Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1474:1470]));
  assign Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1764:1760]));
  assign Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_972_nl = Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_958_nl
      + Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_972_nl = nl_Accum2_acc_972_nl[8:0];
  assign nl_Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3214:3210]));
  assign Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3504:3500]));
  assign Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2054:2050]));
  assign Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2344:2340]));
  assign Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2634:2630]));
  assign Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2924:2920]));
  assign Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3794:3790]));
  assign Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4084:4080]));
  assign Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_971_nl = Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_971_nl = nl_Accum2_acc_971_nl[8:0];
  assign nl_Accum2_acc_68_psp_sva_1 = Accum2_acc_972_nl + Accum2_acc_971_nl;
  assign Accum2_acc_68_psp_sva_1 = nl_Accum2_acc_68_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 = (Accum2_acc_69_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[899:895]));
  assign Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1189:1185]));
  assign Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4379:4375]));
  assign Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_973_nl = Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[29:25]);
  assign Accum2_acc_973_nl = nl_Accum2_acc_973_nl[8:0];
  assign nl_Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[29:25]));
  assign Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[319:315]));
  assign Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[609:605]));
  assign Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1479:1475]));
  assign Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1769:1765]));
  assign Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_987_nl = Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_973_nl
      + Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_987_nl = nl_Accum2_acc_987_nl[8:0];
  assign nl_Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3219:3215]));
  assign Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3509:3505]));
  assign Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2059:2055]));
  assign Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2349:2345]));
  assign Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2639:2635]));
  assign Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2929:2925]));
  assign Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3799:3795]));
  assign Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4089:4085]));
  assign Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_986_nl = Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_986_nl = nl_Accum2_acc_986_nl[8:0];
  assign nl_Accum2_acc_69_psp_sva_1 = Accum2_acc_987_nl + Accum2_acc_986_nl;
  assign Accum2_acc_69_psp_sva_1 = nl_Accum2_acc_69_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 = (Accum2_acc_70_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[904:900]));
  assign Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1194:1190]));
  assign Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4384:4380]));
  assign Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_988_nl = Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[34:30]);
  assign Accum2_acc_988_nl = nl_Accum2_acc_988_nl[8:0];
  assign nl_Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[34:30]));
  assign Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[324:320]));
  assign Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[614:610]));
  assign Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1484:1480]));
  assign Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1774:1770]));
  assign Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1002_nl = Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_988_nl
      + Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1002_nl = nl_Accum2_acc_1002_nl[8:0];
  assign nl_Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3224:3220]));
  assign Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3514:3510]));
  assign Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2064:2060]));
  assign Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2354:2350]));
  assign Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2644:2640]));
  assign Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2934:2930]));
  assign Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3804:3800]));
  assign Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4094:4090]));
  assign Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1001_nl = Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1001_nl = nl_Accum2_acc_1001_nl[8:0];
  assign nl_Accum2_acc_70_psp_sva_1 = Accum2_acc_1002_nl + Accum2_acc_1001_nl;
  assign Accum2_acc_70_psp_sva_1 = nl_Accum2_acc_70_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 = (Accum2_acc_71_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[909:905]));
  assign Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1199:1195]));
  assign Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4389:4385]));
  assign Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1003_nl = Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[39:35]);
  assign Accum2_acc_1003_nl = nl_Accum2_acc_1003_nl[8:0];
  assign nl_Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[39:35]));
  assign Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[329:325]));
  assign Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[619:615]));
  assign Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1489:1485]));
  assign Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1779:1775]));
  assign Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1017_nl = Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_1003_nl
      + Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1017_nl = nl_Accum2_acc_1017_nl[8:0];
  assign nl_Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3229:3225]));
  assign Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3519:3515]));
  assign Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2069:2065]));
  assign Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2359:2355]));
  assign Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2649:2645]));
  assign Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2939:2935]));
  assign Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3809:3805]));
  assign Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4099:4095]));
  assign Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1016_nl = Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1016_nl = nl_Accum2_acc_1016_nl[8:0];
  assign nl_Accum2_acc_71_psp_sva_1 = Accum2_acc_1017_nl + Accum2_acc_1016_nl;
  assign Accum2_acc_71_psp_sva_1 = nl_Accum2_acc_71_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 = (Accum2_acc_72_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[914:910]));
  assign Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1204:1200]));
  assign Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4394:4390]));
  assign Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1018_nl = Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[44:40]);
  assign Accum2_acc_1018_nl = nl_Accum2_acc_1018_nl[8:0];
  assign nl_Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[44:40]));
  assign Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[334:330]));
  assign Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[624:620]));
  assign Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1494:1490]));
  assign Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1784:1780]));
  assign Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1032_nl = Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Accum2_acc_1018_nl
      + Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1032_nl = nl_Accum2_acc_1032_nl[8:0];
  assign nl_Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3234:3230]));
  assign Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3524:3520]));
  assign Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2074:2070]));
  assign Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2364:2360]));
  assign Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2654:2650]));
  assign Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2944:2940]));
  assign Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3814:3810]));
  assign Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4104:4100]));
  assign Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1031_nl = Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1031_nl = nl_Accum2_acc_1031_nl[8:0];
  assign nl_Accum2_acc_72_psp_sva_1 = Accum2_acc_1032_nl + Accum2_acc_1031_nl;
  assign Accum2_acc_72_psp_sva_1 = nl_Accum2_acc_72_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 = (Accum2_acc_73_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[919:915]));
  assign Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1209:1205]));
  assign Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4399:4395]));
  assign Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1033_nl = Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[49:45]);
  assign Accum2_acc_1033_nl = nl_Accum2_acc_1033_nl[8:0];
  assign nl_Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[49:45]));
  assign Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[339:335]));
  assign Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[629:625]));
  assign Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1499:1495]));
  assign Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1789:1785]));
  assign Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1047_nl = Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1033_nl + Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1047_nl = nl_Accum2_acc_1047_nl[8:0];
  assign nl_Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3239:3235]));
  assign Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3529:3525]));
  assign Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2079:2075]));
  assign Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2369:2365]));
  assign Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2659:2655]));
  assign Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2949:2945]));
  assign Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3819:3815]));
  assign Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4109:4105]));
  assign Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1046_nl = Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1046_nl = nl_Accum2_acc_1046_nl[8:0];
  assign nl_Accum2_acc_73_psp_sva_1 = Accum2_acc_1047_nl + Accum2_acc_1046_nl;
  assign Accum2_acc_73_psp_sva_1 = nl_Accum2_acc_73_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 = (Accum2_acc_74_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[924:920]));
  assign Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1214:1210]));
  assign Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4404:4400]));
  assign Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1048_nl = Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[54:50]);
  assign Accum2_acc_1048_nl = nl_Accum2_acc_1048_nl[8:0];
  assign nl_Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[54:50]));
  assign Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[344:340]));
  assign Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[634:630]));
  assign Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1504:1500]));
  assign Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1794:1790]));
  assign Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1062_nl = Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1048_nl + Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1062_nl = nl_Accum2_acc_1062_nl[8:0];
  assign nl_Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3244:3240]));
  assign Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3534:3530]));
  assign Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2084:2080]));
  assign Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2374:2370]));
  assign Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2664:2660]));
  assign Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2954:2950]));
  assign Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3824:3820]));
  assign Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4114:4110]));
  assign Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1061_nl = Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1061_nl = nl_Accum2_acc_1061_nl[8:0];
  assign nl_Accum2_acc_74_psp_sva_1 = Accum2_acc_1062_nl + Accum2_acc_1061_nl;
  assign Accum2_acc_74_psp_sva_1 = nl_Accum2_acc_74_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 = (Accum2_acc_75_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[929:925]));
  assign Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1219:1215]));
  assign Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4409:4405]));
  assign Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1063_nl = Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[59:55]);
  assign Accum2_acc_1063_nl = nl_Accum2_acc_1063_nl[8:0];
  assign nl_Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[59:55]));
  assign Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[349:345]));
  assign Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[639:635]));
  assign Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1509:1505]));
  assign Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1799:1795]));
  assign Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1077_nl = Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1063_nl + Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1077_nl = nl_Accum2_acc_1077_nl[8:0];
  assign nl_Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3249:3245]));
  assign Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3539:3535]));
  assign Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2089:2085]));
  assign Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2379:2375]));
  assign Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2669:2665]));
  assign Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2959:2955]));
  assign Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3829:3825]));
  assign Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4119:4115]));
  assign Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1076_nl = Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1076_nl = nl_Accum2_acc_1076_nl[8:0];
  assign nl_Accum2_acc_75_psp_sva_1 = Accum2_acc_1077_nl + Accum2_acc_1076_nl;
  assign Accum2_acc_75_psp_sva_1 = nl_Accum2_acc_75_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 = (Accum2_acc_76_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[934:930]));
  assign Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1224:1220]));
  assign Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4414:4410]));
  assign Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1078_nl = Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[64:60]);
  assign Accum2_acc_1078_nl = nl_Accum2_acc_1078_nl[8:0];
  assign nl_Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[64:60]));
  assign Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[354:350]));
  assign Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[644:640]));
  assign Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1514:1510]));
  assign Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1804:1800]));
  assign Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1092_nl = Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1078_nl + Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1092_nl = nl_Accum2_acc_1092_nl[8:0];
  assign nl_Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3254:3250]));
  assign Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3544:3540]));
  assign Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2094:2090]));
  assign Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2384:2380]));
  assign Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2674:2670]));
  assign Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2964:2960]));
  assign Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3834:3830]));
  assign Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4124:4120]));
  assign Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1091_nl = Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1091_nl = nl_Accum2_acc_1091_nl[8:0];
  assign nl_Accum2_acc_76_psp_sva_1 = Accum2_acc_1092_nl + Accum2_acc_1091_nl;
  assign Accum2_acc_76_psp_sva_1 = nl_Accum2_acc_76_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 = (Accum2_acc_77_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[939:935]));
  assign Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1229:1225]));
  assign Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4419:4415]));
  assign Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1093_nl = Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[69:65]);
  assign Accum2_acc_1093_nl = nl_Accum2_acc_1093_nl[8:0];
  assign nl_Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[69:65]));
  assign Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[359:355]));
  assign Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[649:645]));
  assign Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1519:1515]));
  assign Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1809:1805]));
  assign Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1107_nl = Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1093_nl + Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1107_nl = nl_Accum2_acc_1107_nl[8:0];
  assign nl_Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3259:3255]));
  assign Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3549:3545]));
  assign Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2099:2095]));
  assign Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2389:2385]));
  assign Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2679:2675]));
  assign Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2969:2965]));
  assign Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3839:3835]));
  assign Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4129:4125]));
  assign Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1106_nl = Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1106_nl = nl_Accum2_acc_1106_nl[8:0];
  assign nl_Accum2_acc_77_psp_sva_1 = Accum2_acc_1107_nl + Accum2_acc_1106_nl;
  assign Accum2_acc_77_psp_sva_1 = nl_Accum2_acc_77_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 = (Accum2_acc_78_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[944:940]));
  assign Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1234:1230]));
  assign Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4424:4420]));
  assign Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1108_nl = Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[74:70]);
  assign Accum2_acc_1108_nl = nl_Accum2_acc_1108_nl[8:0];
  assign nl_Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[74:70]));
  assign Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[364:360]));
  assign Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[654:650]));
  assign Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1524:1520]));
  assign Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1814:1810]));
  assign Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1122_nl = Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1108_nl + Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1122_nl = nl_Accum2_acc_1122_nl[8:0];
  assign nl_Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3264:3260]));
  assign Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3554:3550]));
  assign Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2104:2100]));
  assign Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2394:2390]));
  assign Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2684:2680]));
  assign Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2974:2970]));
  assign Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3844:3840]));
  assign Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4134:4130]));
  assign Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1121_nl = Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1121_nl = nl_Accum2_acc_1121_nl[8:0];
  assign nl_Accum2_acc_78_psp_sva_1 = Accum2_acc_1122_nl + Accum2_acc_1121_nl;
  assign Accum2_acc_78_psp_sva_1 = nl_Accum2_acc_78_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 = (Accum2_acc_79_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[949:945]));
  assign Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1239:1235]));
  assign Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4429:4425]));
  assign Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1123_nl = Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[79:75]);
  assign Accum2_acc_1123_nl = nl_Accum2_acc_1123_nl[8:0];
  assign nl_Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[79:75]));
  assign Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[369:365]));
  assign Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[659:655]));
  assign Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1529:1525]));
  assign Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1819:1815]));
  assign Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1137_nl = Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1123_nl + Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1137_nl = nl_Accum2_acc_1137_nl[8:0];
  assign nl_Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3269:3265]));
  assign Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3559:3555]));
  assign Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2109:2105]));
  assign Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2399:2395]));
  assign Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2689:2685]));
  assign Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2979:2975]));
  assign Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3849:3845]));
  assign Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4139:4135]));
  assign Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1136_nl = Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1136_nl = nl_Accum2_acc_1136_nl[8:0];
  assign nl_Accum2_acc_79_psp_sva_1 = Accum2_acc_1137_nl + Accum2_acc_1136_nl;
  assign Accum2_acc_79_psp_sva_1 = nl_Accum2_acc_79_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 = (Accum2_acc_80_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[954:950]));
  assign Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1244:1240]));
  assign Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4434:4430]));
  assign Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1138_nl = Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[84:80]);
  assign Accum2_acc_1138_nl = nl_Accum2_acc_1138_nl[8:0];
  assign nl_Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[84:80]));
  assign Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[374:370]));
  assign Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[664:660]));
  assign Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1534:1530]));
  assign Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1824:1820]));
  assign Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1152_nl = Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1138_nl + Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1152_nl = nl_Accum2_acc_1152_nl[8:0];
  assign nl_Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3274:3270]));
  assign Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3564:3560]));
  assign Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2114:2110]));
  assign Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2404:2400]));
  assign Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2694:2690]));
  assign Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2984:2980]));
  assign Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3854:3850]));
  assign Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4144:4140]));
  assign Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1151_nl = Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1151_nl = nl_Accum2_acc_1151_nl[8:0];
  assign nl_Accum2_acc_80_psp_sva_1 = Accum2_acc_1152_nl + Accum2_acc_1151_nl;
  assign Accum2_acc_80_psp_sva_1 = nl_Accum2_acc_80_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 = (Accum2_acc_81_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[959:955]));
  assign Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1249:1245]));
  assign Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4439:4435]));
  assign Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1153_nl = Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[89:85]);
  assign Accum2_acc_1153_nl = nl_Accum2_acc_1153_nl[8:0];
  assign nl_Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[89:85]));
  assign Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[379:375]));
  assign Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[669:665]));
  assign Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1539:1535]));
  assign Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1829:1825]));
  assign Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1167_nl = Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1153_nl + Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1167_nl = nl_Accum2_acc_1167_nl[8:0];
  assign nl_Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3279:3275]));
  assign Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3569:3565]));
  assign Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2119:2115]));
  assign Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2409:2405]));
  assign Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2699:2695]));
  assign Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2989:2985]));
  assign Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3859:3855]));
  assign Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4149:4145]));
  assign Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1166_nl = Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1166_nl = nl_Accum2_acc_1166_nl[8:0];
  assign nl_Accum2_acc_81_psp_sva_1 = Accum2_acc_1167_nl + Accum2_acc_1166_nl;
  assign Accum2_acc_81_psp_sva_1 = nl_Accum2_acc_81_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 = (Accum2_acc_82_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[964:960]));
  assign Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1254:1250]));
  assign Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4444:4440]));
  assign Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1168_nl = Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[94:90]);
  assign Accum2_acc_1168_nl = nl_Accum2_acc_1168_nl[8:0];
  assign nl_Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[94:90]));
  assign Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[384:380]));
  assign Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[674:670]));
  assign Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1544:1540]));
  assign Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1834:1830]));
  assign Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1182_nl = Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1168_nl + Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1182_nl = nl_Accum2_acc_1182_nl[8:0];
  assign nl_Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3284:3280]));
  assign Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3574:3570]));
  assign Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2124:2120]));
  assign Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2414:2410]));
  assign Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2704:2700]));
  assign Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2994:2990]));
  assign Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3864:3860]));
  assign Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4154:4150]));
  assign Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1181_nl = Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1181_nl = nl_Accum2_acc_1181_nl[8:0];
  assign nl_Accum2_acc_82_psp_sva_1 = Accum2_acc_1182_nl + Accum2_acc_1181_nl;
  assign Accum2_acc_82_psp_sva_1 = nl_Accum2_acc_82_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 = (Accum2_acc_83_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[969:965]));
  assign Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1259:1255]));
  assign Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4449:4445]));
  assign Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1183_nl = Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[99:95]);
  assign Accum2_acc_1183_nl = nl_Accum2_acc_1183_nl[8:0];
  assign nl_Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[99:95]));
  assign Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[389:385]));
  assign Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[679:675]));
  assign Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1549:1545]));
  assign Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1839:1835]));
  assign Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1197_nl = Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1183_nl + Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1197_nl = nl_Accum2_acc_1197_nl[8:0];
  assign nl_Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3289:3285]));
  assign Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3579:3575]));
  assign Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2129:2125]));
  assign Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2419:2415]));
  assign Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2709:2705]));
  assign Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[2999:2995]));
  assign Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3869:3865]));
  assign Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4159:4155]));
  assign Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1196_nl = Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1196_nl = nl_Accum2_acc_1196_nl[8:0];
  assign nl_Accum2_acc_83_psp_sva_1 = Accum2_acc_1197_nl + Accum2_acc_1196_nl;
  assign Accum2_acc_83_psp_sva_1 = nl_Accum2_acc_83_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 = (Accum2_acc_84_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[974:970]));
  assign Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1264:1260]));
  assign Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4454:4450]));
  assign Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1198_nl = Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[104:100]);
  assign Accum2_acc_1198_nl = nl_Accum2_acc_1198_nl[8:0];
  assign nl_Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[104:100]));
  assign Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[394:390]));
  assign Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[684:680]));
  assign Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1554:1550]));
  assign Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1844:1840]));
  assign Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1212_nl = Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1198_nl + Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1212_nl = nl_Accum2_acc_1212_nl[8:0];
  assign nl_Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3294:3290]));
  assign Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3584:3580]));
  assign Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2134:2130]));
  assign Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2424:2420]));
  assign Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2714:2710]));
  assign Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3004:3000]));
  assign Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3874:3870]));
  assign Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4164:4160]));
  assign Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1211_nl = Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1211_nl = nl_Accum2_acc_1211_nl[8:0];
  assign nl_Accum2_acc_84_psp_sva_1 = Accum2_acc_1212_nl + Accum2_acc_1211_nl;
  assign Accum2_acc_84_psp_sva_1 = nl_Accum2_acc_84_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 = (Accum2_acc_85_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[979:975]));
  assign Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1269:1265]));
  assign Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4459:4455]));
  assign Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1213_nl = Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[109:105]);
  assign Accum2_acc_1213_nl = nl_Accum2_acc_1213_nl[8:0];
  assign nl_Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[109:105]));
  assign Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[399:395]));
  assign Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[689:685]));
  assign Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1559:1555]));
  assign Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1849:1845]));
  assign Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1227_nl = Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1213_nl + Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1227_nl = nl_Accum2_acc_1227_nl[8:0];
  assign nl_Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3299:3295]));
  assign Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3589:3585]));
  assign Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2139:2135]));
  assign Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2429:2425]));
  assign Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2719:2715]));
  assign Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3009:3005]));
  assign Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3879:3875]));
  assign Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4169:4165]));
  assign Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1226_nl = Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1226_nl = nl_Accum2_acc_1226_nl[8:0];
  assign nl_Accum2_acc_85_psp_sva_1 = Accum2_acc_1227_nl + Accum2_acc_1226_nl;
  assign Accum2_acc_85_psp_sva_1 = nl_Accum2_acc_85_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 = (Accum2_acc_86_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[984:980]));
  assign Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1274:1270]));
  assign Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4464:4460]));
  assign Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1228_nl = Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[114:110]);
  assign Accum2_acc_1228_nl = nl_Accum2_acc_1228_nl[8:0];
  assign nl_Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[114:110]));
  assign Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[404:400]));
  assign Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[694:690]));
  assign Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1564:1560]));
  assign Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1854:1850]));
  assign Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1242_nl = Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1228_nl + Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1242_nl = nl_Accum2_acc_1242_nl[8:0];
  assign nl_Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3304:3300]));
  assign Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3594:3590]));
  assign Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2144:2140]));
  assign Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2434:2430]));
  assign Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2724:2720]));
  assign Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3014:3010]));
  assign Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3884:3880]));
  assign Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4174:4170]));
  assign Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1241_nl = Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1241_nl = nl_Accum2_acc_1241_nl[8:0];
  assign nl_Accum2_acc_86_psp_sva_1 = Accum2_acc_1242_nl + Accum2_acc_1241_nl;
  assign Accum2_acc_86_psp_sva_1 = nl_Accum2_acc_86_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 = (Accum2_acc_87_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[989:985]));
  assign Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1279:1275]));
  assign Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4469:4465]));
  assign Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1243_nl = Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[119:115]);
  assign Accum2_acc_1243_nl = nl_Accum2_acc_1243_nl[8:0];
  assign nl_Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[119:115]));
  assign Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[409:405]));
  assign Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[699:695]));
  assign Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1569:1565]));
  assign Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1859:1855]));
  assign Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1257_nl = Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1243_nl + Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1257_nl = nl_Accum2_acc_1257_nl[8:0];
  assign nl_Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3309:3305]));
  assign Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3599:3595]));
  assign Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2149:2145]));
  assign Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2439:2435]));
  assign Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2729:2725]));
  assign Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3019:3015]));
  assign Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3889:3885]));
  assign Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4179:4175]));
  assign Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1256_nl = Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1256_nl = nl_Accum2_acc_1256_nl[8:0];
  assign nl_Accum2_acc_87_psp_sva_1 = Accum2_acc_1257_nl + Accum2_acc_1256_nl;
  assign Accum2_acc_87_psp_sva_1 = nl_Accum2_acc_87_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 = (Accum2_acc_88_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[994:990]));
  assign Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1284:1280]));
  assign Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4474:4470]));
  assign Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1258_nl = Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[124:120]);
  assign Accum2_acc_1258_nl = nl_Accum2_acc_1258_nl[8:0];
  assign nl_Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[124:120]));
  assign Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[414:410]));
  assign Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[704:700]));
  assign Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1574:1570]));
  assign Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1864:1860]));
  assign Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1272_nl = Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1258_nl + Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1272_nl = nl_Accum2_acc_1272_nl[8:0];
  assign nl_Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3314:3310]));
  assign Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3604:3600]));
  assign Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2154:2150]));
  assign Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2444:2440]));
  assign Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2734:2730]));
  assign Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3024:3020]));
  assign Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3894:3890]));
  assign Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4184:4180]));
  assign Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1271_nl = Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1271_nl = nl_Accum2_acc_1271_nl[8:0];
  assign nl_Accum2_acc_88_psp_sva_1 = Accum2_acc_1272_nl + Accum2_acc_1271_nl;
  assign Accum2_acc_88_psp_sva_1 = nl_Accum2_acc_88_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 = (Accum2_acc_89_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[999:995]));
  assign Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1289:1285]));
  assign Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4479:4475]));
  assign Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1273_nl = Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[129:125]);
  assign Accum2_acc_1273_nl = nl_Accum2_acc_1273_nl[8:0];
  assign nl_Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[129:125]));
  assign Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[419:415]));
  assign Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[709:705]));
  assign Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1579:1575]));
  assign Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1869:1865]));
  assign Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1287_nl = Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1273_nl + Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1287_nl = nl_Accum2_acc_1287_nl[8:0];
  assign nl_Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3319:3315]));
  assign Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3609:3605]));
  assign Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2159:2155]));
  assign Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2449:2445]));
  assign Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2739:2735]));
  assign Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3029:3025]));
  assign Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3899:3895]));
  assign Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4189:4185]));
  assign Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1286_nl = Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1286_nl = nl_Accum2_acc_1286_nl[8:0];
  assign nl_Accum2_acc_89_psp_sva_1 = Accum2_acc_1287_nl + Accum2_acc_1286_nl;
  assign Accum2_acc_89_psp_sva_1 = nl_Accum2_acc_89_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 = (Accum2_acc_90_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1004:1000]));
  assign Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1294:1290]));
  assign Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4484:4480]));
  assign Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1288_nl = Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[134:130]);
  assign Accum2_acc_1288_nl = nl_Accum2_acc_1288_nl[8:0];
  assign nl_Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[134:130]));
  assign Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[424:420]));
  assign Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[714:710]));
  assign Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1584:1580]));
  assign Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1874:1870]));
  assign Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1302_nl = Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1288_nl + Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1302_nl = nl_Accum2_acc_1302_nl[8:0];
  assign nl_Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3324:3320]));
  assign Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3614:3610]));
  assign Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2164:2160]));
  assign Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2454:2450]));
  assign Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2744:2740]));
  assign Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3034:3030]));
  assign Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3904:3900]));
  assign Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4194:4190]));
  assign Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1301_nl = Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1301_nl = nl_Accum2_acc_1301_nl[8:0];
  assign nl_Accum2_acc_90_psp_sva_1 = Accum2_acc_1302_nl + Accum2_acc_1301_nl;
  assign Accum2_acc_90_psp_sva_1 = nl_Accum2_acc_90_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 = (Accum2_acc_91_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1009:1005]));
  assign Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1299:1295]));
  assign Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4489:4485]));
  assign Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1303_nl = Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[139:135]);
  assign Accum2_acc_1303_nl = nl_Accum2_acc_1303_nl[8:0];
  assign nl_Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[139:135]));
  assign Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[429:425]));
  assign Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[719:715]));
  assign Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1589:1585]));
  assign Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1879:1875]));
  assign Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1317_nl = Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1303_nl + Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1317_nl = nl_Accum2_acc_1317_nl[8:0];
  assign nl_Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3329:3325]));
  assign Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3619:3615]));
  assign Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2169:2165]));
  assign Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2459:2455]));
  assign Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2749:2745]));
  assign Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3039:3035]));
  assign Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3909:3905]));
  assign Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4199:4195]));
  assign Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1316_nl = Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1316_nl = nl_Accum2_acc_1316_nl[8:0];
  assign nl_Accum2_acc_91_psp_sva_1 = Accum2_acc_1317_nl + Accum2_acc_1316_nl;
  assign Accum2_acc_91_psp_sva_1 = nl_Accum2_acc_91_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 = (Accum2_acc_92_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1014:1010]));
  assign Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1304:1300]));
  assign Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4494:4490]));
  assign Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1318_nl = Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[144:140]);
  assign Accum2_acc_1318_nl = nl_Accum2_acc_1318_nl[8:0];
  assign nl_Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[144:140]));
  assign Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[434:430]));
  assign Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[724:720]));
  assign Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1594:1590]));
  assign Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1884:1880]));
  assign Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1332_nl = Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1318_nl + Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1332_nl = nl_Accum2_acc_1332_nl[8:0];
  assign nl_Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3334:3330]));
  assign Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3624:3620]));
  assign Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2174:2170]));
  assign Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2464:2460]));
  assign Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2754:2750]));
  assign Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3044:3040]));
  assign Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3914:3910]));
  assign Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4204:4200]));
  assign Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1331_nl = Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1331_nl = nl_Accum2_acc_1331_nl[8:0];
  assign nl_Accum2_acc_92_psp_sva_1 = Accum2_acc_1332_nl + Accum2_acc_1331_nl;
  assign Accum2_acc_92_psp_sva_1 = nl_Accum2_acc_92_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 = (Accum2_acc_93_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1019:1015]));
  assign Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1309:1305]));
  assign Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4499:4495]));
  assign Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1333_nl = Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[149:145]);
  assign Accum2_acc_1333_nl = nl_Accum2_acc_1333_nl[8:0];
  assign nl_Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[149:145]));
  assign Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[439:435]));
  assign Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[729:725]));
  assign Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1599:1595]));
  assign Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1889:1885]));
  assign Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1347_nl = Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1333_nl + Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1347_nl = nl_Accum2_acc_1347_nl[8:0];
  assign nl_Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3339:3335]));
  assign Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3629:3625]));
  assign Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2179:2175]));
  assign Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2469:2465]));
  assign Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2759:2755]));
  assign Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3049:3045]));
  assign Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3919:3915]));
  assign Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4209:4205]));
  assign Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1346_nl = Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1346_nl = nl_Accum2_acc_1346_nl[8:0];
  assign nl_Accum2_acc_93_psp_sva_1 = Accum2_acc_1347_nl + Accum2_acc_1346_nl;
  assign Accum2_acc_93_psp_sva_1 = nl_Accum2_acc_93_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 = (Accum2_acc_94_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1024:1020]));
  assign Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1314:1310]));
  assign Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4504:4500]));
  assign Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1348_nl = Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[154:150]);
  assign Accum2_acc_1348_nl = nl_Accum2_acc_1348_nl[8:0];
  assign nl_Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[154:150]));
  assign Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[444:440]));
  assign Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[734:730]));
  assign Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1604:1600]));
  assign Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1894:1890]));
  assign Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1362_nl = Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1348_nl + Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1362_nl = nl_Accum2_acc_1362_nl[8:0];
  assign nl_Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3344:3340]));
  assign Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3634:3630]));
  assign Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2184:2180]));
  assign Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2474:2470]));
  assign Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2764:2760]));
  assign Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3054:3050]));
  assign Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3924:3920]));
  assign Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4214:4210]));
  assign Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1361_nl = Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1361_nl = nl_Accum2_acc_1361_nl[8:0];
  assign nl_Accum2_acc_94_psp_sva_1 = Accum2_acc_1362_nl + Accum2_acc_1361_nl;
  assign Accum2_acc_94_psp_sva_1 = nl_Accum2_acc_94_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 = (Accum2_acc_95_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1029:1025]));
  assign Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1319:1315]));
  assign Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4509:4505]));
  assign Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1363_nl = Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[159:155]);
  assign Accum2_acc_1363_nl = nl_Accum2_acc_1363_nl[8:0];
  assign nl_Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[159:155]));
  assign Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[449:445]));
  assign Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[739:735]));
  assign Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1609:1605]));
  assign Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1899:1895]));
  assign Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1377_nl = Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1363_nl + Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1377_nl = nl_Accum2_acc_1377_nl[8:0];
  assign nl_Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3349:3345]));
  assign Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3639:3635]));
  assign Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2189:2185]));
  assign Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2479:2475]));
  assign Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2769:2765]));
  assign Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3059:3055]));
  assign Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3929:3925]));
  assign Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4219:4215]));
  assign Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1376_nl = Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1376_nl = nl_Accum2_acc_1376_nl[8:0];
  assign nl_Accum2_acc_95_psp_sva_1 = Accum2_acc_1377_nl + Accum2_acc_1376_nl;
  assign Accum2_acc_95_psp_sva_1 = nl_Accum2_acc_95_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 = (Accum2_acc_96_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1034:1030]));
  assign Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1324:1320]));
  assign Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4514:4510]));
  assign Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1378_nl = Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[164:160]);
  assign Accum2_acc_1378_nl = nl_Accum2_acc_1378_nl[8:0];
  assign nl_Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[164:160]));
  assign Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[454:450]));
  assign Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[744:740]));
  assign Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1614:1610]));
  assign Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1904:1900]));
  assign Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1392_nl = Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1378_nl + Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1392_nl = nl_Accum2_acc_1392_nl[8:0];
  assign nl_Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3354:3350]));
  assign Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3644:3640]));
  assign Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2194:2190]));
  assign Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2484:2480]));
  assign Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2774:2770]));
  assign Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3064:3060]));
  assign Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3934:3930]));
  assign Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4224:4220]));
  assign Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1391_nl = Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1391_nl = nl_Accum2_acc_1391_nl[8:0];
  assign nl_Accum2_acc_96_psp_sva_1 = Accum2_acc_1392_nl + Accum2_acc_1391_nl;
  assign Accum2_acc_96_psp_sva_1 = nl_Accum2_acc_96_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 = (Accum2_acc_97_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1039:1035]));
  assign Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1329:1325]));
  assign Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4519:4515]));
  assign Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1393_nl = Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[169:165]);
  assign Accum2_acc_1393_nl = nl_Accum2_acc_1393_nl[8:0];
  assign nl_Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[169:165]));
  assign Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[459:455]));
  assign Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[749:745]));
  assign Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1619:1615]));
  assign Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1909:1905]));
  assign Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1407_nl = Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1393_nl + Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1407_nl = nl_Accum2_acc_1407_nl[8:0];
  assign nl_Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3359:3355]));
  assign Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3649:3645]));
  assign Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2199:2195]));
  assign Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2489:2485]));
  assign Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2779:2775]));
  assign Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3069:3065]));
  assign Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3939:3935]));
  assign Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4229:4225]));
  assign Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1406_nl = Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1406_nl = nl_Accum2_acc_1406_nl[8:0];
  assign nl_Accum2_acc_97_psp_sva_1 = Accum2_acc_1407_nl + Accum2_acc_1406_nl;
  assign Accum2_acc_97_psp_sva_1 = nl_Accum2_acc_97_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 = (Accum2_acc_98_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1044:1040]));
  assign Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1334:1330]));
  assign Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4524:4520]));
  assign Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1408_nl = Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[174:170]);
  assign Accum2_acc_1408_nl = nl_Accum2_acc_1408_nl[8:0];
  assign nl_Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[174:170]));
  assign Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[464:460]));
  assign Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[754:750]));
  assign Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1624:1620]));
  assign Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1914:1910]));
  assign Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1422_nl = Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1408_nl + Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1422_nl = nl_Accum2_acc_1422_nl[8:0];
  assign nl_Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3364:3360]));
  assign Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3654:3650]));
  assign Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2204:2200]));
  assign Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2494:2490]));
  assign Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2784:2780]));
  assign Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3074:3070]));
  assign Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3944:3940]));
  assign Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4234:4230]));
  assign Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1421_nl = Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1421_nl = nl_Accum2_acc_1421_nl[8:0];
  assign nl_Accum2_acc_98_psp_sva_1 = Accum2_acc_1422_nl + Accum2_acc_1421_nl;
  assign Accum2_acc_98_psp_sva_1 = nl_Accum2_acc_98_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 = (Accum2_acc_99_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1049:1045]));
  assign Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1339:1335]));
  assign Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4529:4525]));
  assign Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1423_nl = Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[179:175]);
  assign Accum2_acc_1423_nl = nl_Accum2_acc_1423_nl[8:0];
  assign nl_Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[179:175]));
  assign Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[469:465]));
  assign Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[759:755]));
  assign Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1629:1625]));
  assign Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1919:1915]));
  assign Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1437_nl = Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1423_nl + Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1437_nl = nl_Accum2_acc_1437_nl[8:0];
  assign nl_Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3369:3365]));
  assign Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3659:3655]));
  assign Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2209:2205]));
  assign Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2499:2495]));
  assign Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2789:2785]));
  assign Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3079:3075]));
  assign Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3949:3945]));
  assign Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4239:4235]));
  assign Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1436_nl = Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1436_nl = nl_Accum2_acc_1436_nl[8:0];
  assign nl_Accum2_acc_99_psp_sva_1 = Accum2_acc_1437_nl + Accum2_acc_1436_nl;
  assign Accum2_acc_99_psp_sva_1 = nl_Accum2_acc_99_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 = (Accum2_acc_100_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1054:1050]));
  assign Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1344:1340]));
  assign Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4534:4530]));
  assign Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1438_nl = Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[184:180]);
  assign Accum2_acc_1438_nl = nl_Accum2_acc_1438_nl[8:0];
  assign nl_Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[184:180]));
  assign Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[474:470]));
  assign Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[764:760]));
  assign Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1634:1630]));
  assign Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1924:1920]));
  assign Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1452_nl = Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1438_nl + Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1452_nl = nl_Accum2_acc_1452_nl[8:0];
  assign nl_Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3374:3370]));
  assign Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3664:3660]));
  assign Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2214:2210]));
  assign Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2504:2500]));
  assign Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2794:2790]));
  assign Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3084:3080]));
  assign Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3954:3950]));
  assign Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4244:4240]));
  assign Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1451_nl = Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1451_nl = nl_Accum2_acc_1451_nl[8:0];
  assign nl_Accum2_acc_100_psp_sva_1 = Accum2_acc_1452_nl + Accum2_acc_1451_nl;
  assign Accum2_acc_100_psp_sva_1 = nl_Accum2_acc_100_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 = (Accum2_acc_101_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1059:1055]));
  assign Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1349:1345]));
  assign Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4539:4535]));
  assign Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1453_nl = Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[189:185]);
  assign Accum2_acc_1453_nl = nl_Accum2_acc_1453_nl[8:0];
  assign nl_Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[189:185]));
  assign Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[479:475]));
  assign Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[769:765]));
  assign Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1639:1635]));
  assign Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1929:1925]));
  assign Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1467_nl = Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1453_nl + Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1467_nl = nl_Accum2_acc_1467_nl[8:0];
  assign nl_Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3379:3375]));
  assign Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3669:3665]));
  assign Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2219:2215]));
  assign Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2509:2505]));
  assign Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2799:2795]));
  assign Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3089:3085]));
  assign Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3959:3955]));
  assign Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4249:4245]));
  assign Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1466_nl = Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1466_nl = nl_Accum2_acc_1466_nl[8:0];
  assign nl_Accum2_acc_101_psp_sva_1 = Accum2_acc_1467_nl + Accum2_acc_1466_nl;
  assign Accum2_acc_101_psp_sva_1 = nl_Accum2_acc_101_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 = (Accum2_acc_102_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1064:1060]));
  assign Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1354:1350]));
  assign Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4544:4540]));
  assign Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1468_nl = Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[194:190]);
  assign Accum2_acc_1468_nl = nl_Accum2_acc_1468_nl[8:0];
  assign nl_Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[194:190]));
  assign Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[484:480]));
  assign Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[774:770]));
  assign Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1644:1640]));
  assign Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1934:1930]));
  assign Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1482_nl = Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1468_nl + Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1482_nl = nl_Accum2_acc_1482_nl[8:0];
  assign nl_Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3384:3380]));
  assign Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3674:3670]));
  assign Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2224:2220]));
  assign Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2514:2510]));
  assign Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2804:2800]));
  assign Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3094:3090]));
  assign Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3964:3960]));
  assign Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4254:4250]));
  assign Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1481_nl = Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1481_nl = nl_Accum2_acc_1481_nl[8:0];
  assign nl_Accum2_acc_102_psp_sva_1 = Accum2_acc_1482_nl + Accum2_acc_1481_nl;
  assign Accum2_acc_102_psp_sva_1 = nl_Accum2_acc_102_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 = (Accum2_acc_103_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1069:1065]));
  assign Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1359:1355]));
  assign Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4549:4545]));
  assign Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1483_nl = Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[199:195]);
  assign Accum2_acc_1483_nl = nl_Accum2_acc_1483_nl[8:0];
  assign nl_Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[199:195]));
  assign Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[489:485]));
  assign Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[779:775]));
  assign Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1649:1645]));
  assign Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1939:1935]));
  assign Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1497_nl = Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1483_nl + Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1497_nl = nl_Accum2_acc_1497_nl[8:0];
  assign nl_Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3389:3385]));
  assign Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3679:3675]));
  assign Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2229:2225]));
  assign Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2519:2515]));
  assign Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2809:2805]));
  assign Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3099:3095]));
  assign Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3969:3965]));
  assign Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4259:4255]));
  assign Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1496_nl = Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1496_nl = nl_Accum2_acc_1496_nl[8:0];
  assign nl_Accum2_acc_103_psp_sva_1 = Accum2_acc_1497_nl + Accum2_acc_1496_nl;
  assign Accum2_acc_103_psp_sva_1 = nl_Accum2_acc_103_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 = (Accum2_acc_104_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1074:1070]));
  assign Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1364:1360]));
  assign Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4554:4550]));
  assign Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1498_nl = Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[204:200]);
  assign Accum2_acc_1498_nl = nl_Accum2_acc_1498_nl[8:0];
  assign nl_Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[204:200]));
  assign Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[494:490]));
  assign Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[784:780]));
  assign Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1654:1650]));
  assign Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1944:1940]));
  assign Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1512_nl = Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1498_nl + Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1512_nl = nl_Accum2_acc_1512_nl[8:0];
  assign nl_Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3394:3390]));
  assign Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3684:3680]));
  assign Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2234:2230]));
  assign Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2524:2520]));
  assign Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2814:2810]));
  assign Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3104:3100]));
  assign Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3974:3970]));
  assign Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4264:4260]));
  assign Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1511_nl = Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1511_nl = nl_Accum2_acc_1511_nl[8:0];
  assign nl_Accum2_acc_104_psp_sva_1 = Accum2_acc_1512_nl + Accum2_acc_1511_nl;
  assign Accum2_acc_104_psp_sva_1 = nl_Accum2_acc_104_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 = (Accum2_acc_105_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1079:1075]));
  assign Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1369:1365]));
  assign Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4559:4555]));
  assign Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1513_nl = Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[209:205]);
  assign Accum2_acc_1513_nl = nl_Accum2_acc_1513_nl[8:0];
  assign nl_Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[209:205]));
  assign Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[499:495]));
  assign Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[789:785]));
  assign Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1659:1655]));
  assign Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1949:1945]));
  assign Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1527_nl = Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1513_nl + Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1527_nl = nl_Accum2_acc_1527_nl[8:0];
  assign nl_Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3399:3395]));
  assign Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3689:3685]));
  assign Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2239:2235]));
  assign Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2529:2525]));
  assign Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2819:2815]));
  assign Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3109:3105]));
  assign Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3979:3975]));
  assign Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4269:4265]));
  assign Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1526_nl = Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1526_nl = nl_Accum2_acc_1526_nl[8:0];
  assign nl_Accum2_acc_105_psp_sva_1 = Accum2_acc_1527_nl + Accum2_acc_1526_nl;
  assign Accum2_acc_105_psp_sva_1 = nl_Accum2_acc_105_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 = (Accum2_acc_106_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1084:1080]));
  assign Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1374:1370]));
  assign Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4564:4560]));
  assign Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1528_nl = Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[214:210]);
  assign Accum2_acc_1528_nl = nl_Accum2_acc_1528_nl[8:0];
  assign nl_Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[214:210]));
  assign Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[504:500]));
  assign Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[794:790]));
  assign Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1664:1660]));
  assign Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1954:1950]));
  assign Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1542_nl = Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1528_nl + Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1542_nl = nl_Accum2_acc_1542_nl[8:0];
  assign nl_Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3404:3400]));
  assign Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3694:3690]));
  assign Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2244:2240]));
  assign Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2534:2530]));
  assign Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2824:2820]));
  assign Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3114:3110]));
  assign Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3984:3980]));
  assign Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4274:4270]));
  assign Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1541_nl = Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1541_nl = nl_Accum2_acc_1541_nl[8:0];
  assign nl_Accum2_acc_106_psp_sva_1 = Accum2_acc_1542_nl + Accum2_acc_1541_nl;
  assign Accum2_acc_106_psp_sva_1 = nl_Accum2_acc_106_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 = (Accum2_acc_107_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1089:1085]));
  assign Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1379:1375]));
  assign Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4569:4565]));
  assign Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1543_nl = Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[219:215]);
  assign Accum2_acc_1543_nl = nl_Accum2_acc_1543_nl[8:0];
  assign nl_Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[219:215]));
  assign Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[509:505]));
  assign Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[799:795]));
  assign Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1669:1665]));
  assign Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1959:1955]));
  assign Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1557_nl = Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1543_nl + Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1557_nl = nl_Accum2_acc_1557_nl[8:0];
  assign nl_Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3409:3405]));
  assign Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3699:3695]));
  assign Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2249:2245]));
  assign Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2539:2535]));
  assign Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2829:2825]));
  assign Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3119:3115]));
  assign Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3989:3985]));
  assign Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4279:4275]));
  assign Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1556_nl = Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1556_nl = nl_Accum2_acc_1556_nl[8:0];
  assign nl_Accum2_acc_107_psp_sva_1 = Accum2_acc_1557_nl + Accum2_acc_1556_nl;
  assign Accum2_acc_107_psp_sva_1 = nl_Accum2_acc_107_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 = (Accum2_acc_108_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1094:1090]));
  assign Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1384:1380]));
  assign Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4574:4570]));
  assign Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1558_nl = Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[224:220]);
  assign Accum2_acc_1558_nl = nl_Accum2_acc_1558_nl[8:0];
  assign nl_Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[224:220]));
  assign Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[514:510]));
  assign Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[804:800]));
  assign Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1674:1670]));
  assign Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1964:1960]));
  assign Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1572_nl = Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1558_nl + Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1572_nl = nl_Accum2_acc_1572_nl[8:0];
  assign nl_Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3414:3410]));
  assign Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3704:3700]));
  assign Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2254:2250]));
  assign Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2544:2540]));
  assign Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2834:2830]));
  assign Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3124:3120]));
  assign Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3994:3990]));
  assign Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4284:4280]));
  assign Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1571_nl = Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1571_nl = nl_Accum2_acc_1571_nl[8:0];
  assign nl_Accum2_acc_108_psp_sva_1 = Accum2_acc_1572_nl + Accum2_acc_1571_nl;
  assign Accum2_acc_108_psp_sva_1 = nl_Accum2_acc_108_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 = (Accum2_acc_109_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1099:1095]));
  assign Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1389:1385]));
  assign Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4579:4575]));
  assign Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1573_nl = Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[229:225]);
  assign Accum2_acc_1573_nl = nl_Accum2_acc_1573_nl[8:0];
  assign nl_Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[229:225]));
  assign Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[519:515]));
  assign Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[809:805]));
  assign Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1679:1675]));
  assign Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1969:1965]));
  assign Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1587_nl = Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1573_nl + Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1587_nl = nl_Accum2_acc_1587_nl[8:0];
  assign nl_Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3419:3415]));
  assign Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3709:3705]));
  assign Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2259:2255]));
  assign Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2549:2545]));
  assign Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2839:2835]));
  assign Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3129:3125]));
  assign Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[3999:3995]));
  assign Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4289:4285]));
  assign Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1586_nl = Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1586_nl = nl_Accum2_acc_1586_nl[8:0];
  assign nl_Accum2_acc_109_psp_sva_1 = Accum2_acc_1587_nl + Accum2_acc_1586_nl;
  assign Accum2_acc_109_psp_sva_1 = nl_Accum2_acc_109_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 = (Accum2_acc_110_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1104:1100]));
  assign Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1394:1390]));
  assign Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4584:4580]));
  assign Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1588_nl = Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[234:230]);
  assign Accum2_acc_1588_nl = nl_Accum2_acc_1588_nl[8:0];
  assign nl_Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[234:230]));
  assign Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[524:520]));
  assign Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[814:810]));
  assign Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1684:1680]));
  assign Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1974:1970]));
  assign Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1602_nl = Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1588_nl + Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1602_nl = nl_Accum2_acc_1602_nl[8:0];
  assign nl_Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3424:3420]));
  assign Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3714:3710]));
  assign Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2264:2260]));
  assign Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2554:2550]));
  assign Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2844:2840]));
  assign Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3134:3130]));
  assign Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4004:4000]));
  assign Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4294:4290]));
  assign Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1601_nl = Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1601_nl = nl_Accum2_acc_1601_nl[8:0];
  assign nl_Accum2_acc_110_psp_sva_1 = Accum2_acc_1602_nl + Accum2_acc_1601_nl;
  assign Accum2_acc_110_psp_sva_1 = nl_Accum2_acc_110_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 = (Accum2_acc_111_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1109:1105]));
  assign Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1399:1395]));
  assign Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4589:4585]));
  assign Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1603_nl = Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[239:235]);
  assign Accum2_acc_1603_nl = nl_Accum2_acc_1603_nl[8:0];
  assign nl_Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[239:235]));
  assign Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[529:525]));
  assign Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[819:815]));
  assign Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1689:1685]));
  assign Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1979:1975]));
  assign Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1617_nl = Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1603_nl + Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1617_nl = nl_Accum2_acc_1617_nl[8:0];
  assign nl_Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3429:3425]));
  assign Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3719:3715]));
  assign Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2269:2265]));
  assign Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2559:2555]));
  assign Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2849:2845]));
  assign Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3139:3135]));
  assign Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4009:4005]));
  assign Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4299:4295]));
  assign Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1616_nl = Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1616_nl = nl_Accum2_acc_1616_nl[8:0];
  assign nl_Accum2_acc_111_psp_sva_1 = Accum2_acc_1617_nl + Accum2_acc_1616_nl;
  assign Accum2_acc_111_psp_sva_1 = nl_Accum2_acc_111_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 = (Accum2_acc_112_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1114:1110]));
  assign Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1404:1400]));
  assign Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4594:4590]));
  assign Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1618_nl = Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[244:240]);
  assign Accum2_acc_1618_nl = nl_Accum2_acc_1618_nl[8:0];
  assign nl_Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[244:240]));
  assign Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[534:530]));
  assign Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[824:820]));
  assign Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1694:1690]));
  assign Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1984:1980]));
  assign Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1632_nl = Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1618_nl + Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1632_nl = nl_Accum2_acc_1632_nl[8:0];
  assign nl_Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3434:3430]));
  assign Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3724:3720]));
  assign Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2274:2270]));
  assign Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2564:2560]));
  assign Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2854:2850]));
  assign Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3144:3140]));
  assign Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4014:4010]));
  assign Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4304:4300]));
  assign Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1631_nl = Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1631_nl = nl_Accum2_acc_1631_nl[8:0];
  assign nl_Accum2_acc_112_psp_sva_1 = Accum2_acc_1632_nl + Accum2_acc_1631_nl;
  assign Accum2_acc_112_psp_sva_1 = nl_Accum2_acc_112_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 = (Accum2_acc_113_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1119:1115]));
  assign Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1409:1405]));
  assign Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4599:4595]));
  assign Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1633_nl = Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[249:245]);
  assign Accum2_acc_1633_nl = nl_Accum2_acc_1633_nl[8:0];
  assign nl_Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[249:245]));
  assign Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[539:535]));
  assign Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[829:825]));
  assign Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1699:1695]));
  assign Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1989:1985]));
  assign Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1647_nl = Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1633_nl + Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1647_nl = nl_Accum2_acc_1647_nl[8:0];
  assign nl_Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3439:3435]));
  assign Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3729:3725]));
  assign Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2279:2275]));
  assign Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2569:2565]));
  assign Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2859:2855]));
  assign Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3149:3145]));
  assign Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4019:4015]));
  assign Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4309:4305]));
  assign Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1646_nl = Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1646_nl = nl_Accum2_acc_1646_nl[8:0];
  assign nl_Accum2_acc_113_psp_sva_1 = Accum2_acc_1647_nl + Accum2_acc_1646_nl;
  assign Accum2_acc_113_psp_sva_1 = nl_Accum2_acc_113_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 = (Accum2_acc_114_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1124:1120]));
  assign Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1414:1410]));
  assign Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4604:4600]));
  assign Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1648_nl = Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[254:250]);
  assign Accum2_acc_1648_nl = nl_Accum2_acc_1648_nl[8:0];
  assign nl_Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[254:250]));
  assign Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[544:540]));
  assign Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[834:830]));
  assign Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1704:1700]));
  assign Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1994:1990]));
  assign Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1662_nl = Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1648_nl + Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1662_nl = nl_Accum2_acc_1662_nl[8:0];
  assign nl_Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3444:3440]));
  assign Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3734:3730]));
  assign Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2284:2280]));
  assign Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2574:2570]));
  assign Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2864:2860]));
  assign Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3154:3150]));
  assign Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4024:4020]));
  assign Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4314:4310]));
  assign Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1661_nl = Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1661_nl = nl_Accum2_acc_1661_nl[8:0];
  assign nl_Accum2_acc_114_psp_sva_1 = Accum2_acc_1662_nl + Accum2_acc_1661_nl;
  assign Accum2_acc_114_psp_sva_1 = nl_Accum2_acc_114_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 = (Accum2_acc_115_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1129:1125]));
  assign Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1419:1415]));
  assign Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4609:4605]));
  assign Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1663_nl = Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[259:255]);
  assign Accum2_acc_1663_nl = nl_Accum2_acc_1663_nl[8:0];
  assign nl_Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[259:255]));
  assign Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[549:545]));
  assign Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[839:835]));
  assign Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1709:1705]));
  assign Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1999:1995]));
  assign Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1677_nl = Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1663_nl + Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1677_nl = nl_Accum2_acc_1677_nl[8:0];
  assign nl_Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3449:3445]));
  assign Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3739:3735]));
  assign Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2289:2285]));
  assign Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2579:2575]));
  assign Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2869:2865]));
  assign Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3159:3155]));
  assign Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4029:4025]));
  assign Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4319:4315]));
  assign Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1676_nl = Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1676_nl = nl_Accum2_acc_1676_nl[8:0];
  assign nl_Accum2_acc_115_psp_sva_1 = Accum2_acc_1677_nl + Accum2_acc_1676_nl;
  assign Accum2_acc_115_psp_sva_1 = nl_Accum2_acc_115_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 = (Accum2_acc_116_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1134:1130]));
  assign Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1424:1420]));
  assign Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4614:4610]));
  assign Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1678_nl = Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[264:260]);
  assign Accum2_acc_1678_nl = nl_Accum2_acc_1678_nl[8:0];
  assign nl_Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[264:260]));
  assign Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[554:550]));
  assign Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[844:840]));
  assign Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1714:1710]));
  assign Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2004:2000]));
  assign Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1692_nl = Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1678_nl + Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1692_nl = nl_Accum2_acc_1692_nl[8:0];
  assign nl_Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3454:3450]));
  assign Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3744:3740]));
  assign Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2294:2290]));
  assign Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2584:2580]));
  assign Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2874:2870]));
  assign Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3164:3160]));
  assign Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4034:4030]));
  assign Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4324:4320]));
  assign Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1691_nl = Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1691_nl = nl_Accum2_acc_1691_nl[8:0];
  assign nl_Accum2_acc_116_psp_sva_1 = Accum2_acc_1692_nl + Accum2_acc_1691_nl;
  assign Accum2_acc_116_psp_sva_1 = nl_Accum2_acc_116_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 = (Accum2_acc_117_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1139:1135]));
  assign Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1429:1425]));
  assign Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4619:4615]));
  assign Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1693_nl = Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[269:265]);
  assign Accum2_acc_1693_nl = nl_Accum2_acc_1693_nl[8:0];
  assign nl_Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[269:265]));
  assign Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[559:555]));
  assign Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[849:845]));
  assign Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1719:1715]));
  assign Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2009:2005]));
  assign Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1707_nl = Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1693_nl + Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1707_nl = nl_Accum2_acc_1707_nl[8:0];
  assign nl_Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3459:3455]));
  assign Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3749:3745]));
  assign Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2299:2295]));
  assign Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2589:2585]));
  assign Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2879:2875]));
  assign Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3169:3165]));
  assign Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4039:4035]));
  assign Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4329:4325]));
  assign Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1706_nl = Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1706_nl = nl_Accum2_acc_1706_nl[8:0];
  assign nl_Accum2_acc_117_psp_sva_1 = Accum2_acc_1707_nl + Accum2_acc_1706_nl;
  assign Accum2_acc_117_psp_sva_1 = nl_Accum2_acc_117_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 = (Accum2_acc_118_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1144:1140]));
  assign Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1434:1430]));
  assign Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4624:4620]));
  assign Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1708_nl = Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[274:270]);
  assign Accum2_acc_1708_nl = nl_Accum2_acc_1708_nl[8:0];
  assign nl_Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[274:270]));
  assign Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[564:560]));
  assign Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[854:850]));
  assign Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1724:1720]));
  assign Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2014:2010]));
  assign Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1722_nl = Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1708_nl + Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1722_nl = nl_Accum2_acc_1722_nl[8:0];
  assign nl_Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3464:3460]));
  assign Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3754:3750]));
  assign Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2304:2300]));
  assign Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2594:2590]));
  assign Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2884:2880]));
  assign Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3174:3170]));
  assign Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4044:4040]));
  assign Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4334:4330]));
  assign Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1721_nl = Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1721_nl = nl_Accum2_acc_1721_nl[8:0];
  assign nl_Accum2_acc_118_psp_sva_1 = Accum2_acc_1722_nl + Accum2_acc_1721_nl;
  assign Accum2_acc_118_psp_sva_1 = nl_Accum2_acc_118_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 = (Accum2_acc_119_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1149:1145]));
  assign Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1439:1435]));
  assign Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4629:4625]));
  assign Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1723_nl = Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[279:275]);
  assign Accum2_acc_1723_nl = nl_Accum2_acc_1723_nl[8:0];
  assign nl_Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[279:275]));
  assign Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[569:565]));
  assign Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[859:855]));
  assign Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1729:1725]));
  assign Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2019:2015]));
  assign Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1737_nl = Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1723_nl + Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1737_nl = nl_Accum2_acc_1737_nl[8:0];
  assign nl_Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3469:3465]));
  assign Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3759:3755]));
  assign Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2309:2305]));
  assign Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2599:2595]));
  assign Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2889:2885]));
  assign Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3179:3175]));
  assign Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4049:4045]));
  assign Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4339:4335]));
  assign Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1736_nl = Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1736_nl = nl_Accum2_acc_1736_nl[8:0];
  assign nl_Accum2_acc_119_psp_sva_1 = Accum2_acc_1737_nl + Accum2_acc_1736_nl;
  assign Accum2_acc_119_psp_sva_1 = nl_Accum2_acc_119_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 = (Accum2_acc_120_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1154:1150]));
  assign Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1444:1440]));
  assign Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4634:4630]));
  assign Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1738_nl = Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[284:280]);
  assign Accum2_acc_1738_nl = nl_Accum2_acc_1738_nl[8:0];
  assign nl_Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[284:280]));
  assign Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[574:570]));
  assign Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[864:860]));
  assign Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1734:1730]));
  assign Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2024:2020]));
  assign Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1752_nl = Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1738_nl + Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1752_nl = nl_Accum2_acc_1752_nl[8:0];
  assign nl_Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3474:3470]));
  assign Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3764:3760]));
  assign Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2314:2310]));
  assign Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2604:2600]));
  assign Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2894:2890]));
  assign Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3184:3180]));
  assign Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4054:4050]));
  assign Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4344:4340]));
  assign Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1751_nl = Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1751_nl = nl_Accum2_acc_1751_nl[8:0];
  assign nl_Accum2_acc_120_psp_sva_1 = Accum2_acc_1752_nl + Accum2_acc_1751_nl;
  assign Accum2_acc_120_psp_sva_1 = nl_Accum2_acc_120_psp_sva_1[8:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 = (Accum2_acc_121_psp_sva_1[7:4]!=4'b0000);
  assign nl_Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1159:1155]));
  assign Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1449:1445]));
  assign Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4639:4635]));
  assign Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1753_nl = Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_9(b2_rsci_idat[289:285]);
  assign Accum2_acc_1753_nl = nl_Accum2_acc_1753_nl[8:0];
  assign nl_Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[289:285]));
  assign Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[579:575]));
  assign Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[869:865]));
  assign Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1739:1735]));
  assign Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2029:2025]));
  assign Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1767_nl = Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Accum2_acc_1753_nl + Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1767_nl = nl_Accum2_acc_1767_nl[8:0];
  assign nl_Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3479:3475]));
  assign Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3769:3765]));
  assign Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2319:2315]));
  assign Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2609:2605]));
  assign Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2899:2895]));
  assign Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3189:3185]));
  assign Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4059:4055]));
  assign Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4349:4345]));
  assign Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[8:0];
  assign nl_Accum2_acc_1766_nl = Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl +
      Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl + Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  assign Accum2_acc_1766_nl = nl_Accum2_acc_1766_nl[8:0];
  assign nl_Accum2_acc_121_psp_sva_1 = Accum2_acc_1767_nl + Accum2_acc_1766_nl;
  assign Accum2_acc_121_psp_sva_1 = nl_Accum2_acc_121_psp_sva_1[8:0];
  assign nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[294:290]));
  assign Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[309:305]));
  assign Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[414:410]));
  assign Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[429:425]));
  assign Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[354:350]));
  assign Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[369:365]));
  assign Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[864:860]));
  assign Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[819:815]));
  assign Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[834:830]));
  assign Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[789:785]));
  assign Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[474:470]));
  assign Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[489:485]));
  assign Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[504:500]));
  assign Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[519:515]));
  assign Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[849:845]));
  assign Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[534:530]));
  assign Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[549:545]));
  assign Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[234:230]));
  assign Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[249:245]));
  assign Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[264:260]));
  assign Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[279:275]));
  assign Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[324:320]));
  assign Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[339:335]));
  assign Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[384:380]));
  assign Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[399:395]));
  assign Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[444:440]));
  assign Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[459:455]));
  assign Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_114_nl = conv_s2s_9_13(readslicef_15_9_6(Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum2_1_acc_114_nl = nl_Accum2_1_acc_114_nl[12:0];
  assign nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[624:620]));
  assign Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[579:575]));
  assign Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[684:680]));
  assign Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[639:635]));
  assign Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[804:800]));
  assign Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[759:755]));
  assign Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[774:770]));
  assign Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[729:725]));
  assign Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[744:740]));
  assign Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[699:695]));
  assign Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[714:710]));
  assign Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[669:665]));
  assign Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_174_nl = conv_s2s_5_6(b5_rsci_idat[9:5]) + conv_s2s_5_6(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[8:4]);
  assign Accum2_1_acc_174_nl = nl_Accum2_1_acc_174_nl[5:0];
  assign nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[24:20]));
  assign Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[39:35]));
  assign Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[54:50]));
  assign Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[69:65]));
  assign Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[84:80]));
  assign Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[99:95]));
  assign Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[174:170]));
  assign Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[189:185]));
  assign Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[204:200]));
  assign Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[219:215]));
  assign Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[114:110]));
  assign Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[129:125]));
  assign Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[144:140]));
  assign Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[159:155]));
  assign Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[654:650]));
  assign Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[609:605]));
  assign Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[594:590]));
  assign Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[564:560]));
  assign Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_nl = Accum2_1_acc_114_nl + conv_s2s_9_13(readslicef_15_9_6(Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_10_13({Accum2_1_acc_174_nl , (Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[3:0])})
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_nl = nl_Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_nl[12:0];
  assign Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_itm_12_3_1 = readslicef_13_10_3(Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_nl);
  assign nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[284:280]));
  assign Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[299:295]));
  assign Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[404:400]));
  assign Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[419:415]));
  assign Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[344:340]));
  assign Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[359:355]));
  assign Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[869:865]));
  assign Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[824:820]));
  assign Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[839:835]));
  assign Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[794:790]));
  assign Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[464:460]));
  assign Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[479:475]));
  assign Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[494:490]));
  assign Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[509:505]));
  assign Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[854:850]));
  assign Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[524:520]));
  assign Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[539:535]));
  assign Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[224:220]));
  assign Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[239:235]));
  assign Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[254:250]));
  assign Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[269:265]));
  assign Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[314:310]));
  assign Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[329:325]));
  assign Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[374:370]));
  assign Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[389:385]));
  assign Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[434:430]));
  assign Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[449:445]));
  assign Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_171_nl = conv_s2s_9_13(readslicef_15_9_6(Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum2_1_acc_171_nl = nl_Accum2_1_acc_171_nl[12:0];
  assign nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[629:625]));
  assign Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[584:580]));
  assign Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[689:685]));
  assign Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[644:640]));
  assign Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[809:805]));
  assign Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[764:760]));
  assign Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[779:775]));
  assign Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[734:730]));
  assign Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[749:745]));
  assign Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[704:700]));
  assign Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[719:715]));
  assign Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[674:670]));
  assign Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_175_nl = conv_s2s_5_6(Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[8:4])
      + conv_s2s_5_6(b5_rsci_idat[14:10]);
  assign Accum2_1_acc_175_nl = nl_Accum2_1_acc_175_nl[5:0];
  assign nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_4_9 , layer4_out_conc_4_8_6 , layer4_out_0_3_lpi_1_dfm_1
      , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1
      , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1})) * $signed((w5_rsci_idat[14:10]));
  assign Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[29:25]));
  assign Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[44:40]));
  assign Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[59:55]));
  assign Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[74:70]));
  assign Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[89:85]));
  assign Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[164:160]));
  assign Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[179:175]));
  assign Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[194:190]));
  assign Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[209:205]));
  assign Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[104:100]));
  assign Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[119:115]));
  assign Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[134:130]));
  assign Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[149:145]));
  assign Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[659:655]));
  assign Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[614:610]));
  assign Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[599:595]));
  assign Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[554:550]));
  assign Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_nl = Accum2_1_acc_171_nl + conv_s2s_9_13(readslicef_15_9_6(Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_10_13({Accum2_1_acc_175_nl , (Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[3:0])})
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_nl = nl_Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_nl[12:0];
  assign Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_itm_12_3_1 = readslicef_13_10_3(Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_nl);
  assign nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[289:285]));
  assign Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[304:300]));
  assign Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[409:405]));
  assign Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[424:420]));
  assign Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[349:345]));
  assign Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[364:360]));
  assign Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[859:855]));
  assign Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[814:810]));
  assign Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[829:825]));
  assign Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[784:780]));
  assign Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[469:465]));
  assign Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[484:480]));
  assign Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[499:495]));
  assign Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[514:510]));
  assign Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[844:840]));
  assign Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[529:525]));
  assign Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[544:540]));
  assign Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[229:225]));
  assign Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[244:240]));
  assign Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[259:255]));
  assign Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[274:270]));
  assign Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[319:315]));
  assign Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[334:330]));
  assign Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[379:375]));
  assign Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[394:390]));
  assign Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[439:435]));
  assign Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[454:450]));
  assign Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_nl = conv_s2s_9_13(readslicef_15_9_6(Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum2_1_acc_nl = nl_Accum2_1_acc_nl[12:0];
  assign nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[619:615]));
  assign Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[574:570]));
  assign Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[679:675]));
  assign Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[634:630]));
  assign Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[799:795]));
  assign Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[754:750]));
  assign Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[769:765]));
  assign Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[724:720]));
  assign Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[739:735]));
  assign Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[694:690]));
  assign Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[709:705]));
  assign Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[664:660]));
  assign Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_173_nl = conv_s2s_5_6(b5_rsci_idat[4:0]) + conv_s2s_5_6(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[8:4]);
  assign Accum2_1_acc_173_nl = nl_Accum2_1_acc_173_nl[5:0];
  assign nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[19:15]));
  assign Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[34:30]));
  assign Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[49:45]));
  assign Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[64:60]));
  assign Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[79:75]));
  assign Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[94:90]));
  assign Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[169:165]));
  assign Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[184:180]));
  assign Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[199:195]));
  assign Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[214:210]));
  assign Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[109:105]));
  assign Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[124:120]));
  assign Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[139:135]));
  assign Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[154:150]));
  assign Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[649:645]));
  assign Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[604:600]));
  assign Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[589:585]));
  assign Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[559:555]));
  assign Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_nl = Accum2_1_acc_nl + conv_s2s_9_13(readslicef_15_9_6(Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_10_13({Accum2_1_acc_173_nl , (Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[3:0])})
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_13(readslicef_15_9_6(Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_nl = nl_Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_nl[12:0];
  assign Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_itm_12_3_1 = readslicef_13_10_3(Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_8_6 , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[569:565]));
  assign Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1
      = readslicef_15_9_6(Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign layer4_out_0_3_lpi_1_dfm_1 = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_10_pmx_3_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 & nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_4_9 , layer4_out_conc_4_8_6 , layer4_out_0_3_lpi_1_dfm_1
      , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1
      , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1})) * $signed((w5_rsci_idat[9:5]));
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1
      = readslicef_15_9_6(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_4_9 , layer4_out_conc_4_8_6 , layer4_out_0_3_lpi_1_dfm_1
      , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1
      , layer4_out_0_3_lpi_1_dfm_1 , layer4_out_0_3_lpi_1_dfm_1})) * $signed((w5_rsci_idat[4:0]));
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1
      = readslicef_15_9_6(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_121_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_120_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_119_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_118_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_117_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_116_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_115_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_114_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_113_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_112_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_111_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_110_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_109_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_108_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_107_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_106_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_105_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_104_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_103_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_102_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_101_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_100_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_99_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_98_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_97_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_96_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_95_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_94_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_93_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_92_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_91_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_90_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_89_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_88_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_87_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_86_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_85_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_84_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_83_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_82_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_81_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_80_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_79_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_78_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_77_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_76_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_75_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_74_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_73_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_72_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_71_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_70_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_69_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_68_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_67_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_66_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ Accum2_acc_65_psp_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = conv_s2s_10_11({(~ layer3_out_0_9_1_sva_1) , 1'b1}) + 11'b00000000001;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl[10:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1
      = readslicef_11_1_10(nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_9 = ((Accum2_acc_117_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_117_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_183_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_9 = ((Accum2_acc_114_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_114_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_185_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_9 = ((Accum2_acc_115_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_115_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_187_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_9 = ((Accum2_acc_112_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_112_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_189_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_9 = ((Accum2_acc_113_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_113_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_191_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_9 = ((Accum2_acc_110_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_110_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_193_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_9 = ((Accum2_acc_111_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_111_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_195_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_9 = ((Accum2_acc_108_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_108_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_197_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_9 = ((Accum2_acc_109_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_109_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_199_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_9 = ((Accum2_acc_106_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_106_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_201_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_9 = ((Accum2_acc_107_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_107_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_203_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_9 = ((Accum2_acc_104_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_104_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_205_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_9 = ((Accum2_acc_105_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_105_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_207_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_9 = ((Accum2_acc_102_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_102_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_209_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_9 = ((Accum2_acc_103_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_103_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_211_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_9 = ((Accum2_acc_100_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_100_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_213_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign layer4_out_conc_4_9 = ((layer3_out_0_9_1_sva_1[3]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1)
      & nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((layer3_out_0_9_1_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1);
  assign layer4_out_conc_4_8_6 = MUX_v_3_2_2(3'b000, nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_1_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_9 = ((Accum2_acc_65_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_65_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_215_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_9 = ((Accum2_acc_66_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_66_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_217_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_9 = ((Accum2_acc_67_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_67_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_219_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_9 = ((Accum2_acc_68_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_68_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_221_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_9 = ((Accum2_acc_69_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_69_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_223_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_9 = ((Accum2_acc_70_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_70_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_225_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_9 = ((Accum2_acc_71_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_71_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_227_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_9 = ((Accum2_acc_72_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_72_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_229_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_9 = ((Accum2_acc_73_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_73_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_231_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_9 = ((Accum2_acc_74_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_74_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_233_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_9 = ((Accum2_acc_75_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_75_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_235_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_9 = ((Accum2_acc_76_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_76_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_237_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_9 = ((Accum2_acc_77_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_77_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_239_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_9 = ((Accum2_acc_78_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_78_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_241_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_9 = ((Accum2_acc_79_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_79_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_243_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_9 = ((Accum2_acc_80_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_80_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_245_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_9 = ((Accum2_acc_81_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_81_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_247_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_9 = ((Accum2_acc_82_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_82_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_249_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_9 = ((Accum2_acc_83_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_83_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_251_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_9 = ((Accum2_acc_84_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_84_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_253_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_9 = ((Accum2_acc_85_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_85_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_255_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_9 = ((Accum2_acc_86_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_86_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_257_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_9 = ((Accum2_acc_87_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_87_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_259_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_9 = ((Accum2_acc_88_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_88_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_261_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_9 = ((Accum2_acc_89_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_89_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_263_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_9 = ((Accum2_acc_90_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_90_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_265_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_9 = ((Accum2_acc_91_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_91_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_267_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_9 = ((Accum2_acc_92_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_92_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_269_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_9 = ((Accum2_acc_93_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_93_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_271_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_9 = ((Accum2_acc_94_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_94_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_273_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_9 = ((Accum2_acc_95_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_95_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_275_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_9 = ((Accum2_acc_96_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_96_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_277_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_9 = ((Accum2_acc_97_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_97_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_279_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_9 = ((Accum2_acc_98_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_98_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_281_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_9 = ((Accum2_acc_99_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_99_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_283_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_9 = ((Accum2_acc_120_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_120_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_285_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_9 = ((Accum2_acc_121_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_121_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_287_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_9 = ((Accum2_acc_118_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_118_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_289_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_9 = ((Accum2_acc_119_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_119_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_291_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_9 = ((Accum2_acc_116_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_116_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_293_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_9 = ((Accum2_acc_101_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1) & nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_101_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_295_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_operator_10_5_true_AC_TRN_AC_WRAP_acc_itm_10_1);
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat <= 2'b00;
    end
    else begin
      layer7_out_rsci_idat <= ~(MUX_v_2_2_2(argmax_else_mux_nl, 2'b11, argmax_if_argmax_if_argmax_if_nor_nl));
    end
  end
  assign nl_argmax_else_aif_acc_nl = conv_s2u_10_11(Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_itm_12_3_1)
      - conv_s2u_10_11(Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_itm_12_3_1);
  assign argmax_else_aif_acc_nl = nl_argmax_else_aif_acc_nl[10:0];
  assign nl_argmax_else_acc_nl = conv_s2u_10_11(Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_itm_12_3_1)
      - conv_s2u_10_11(Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_itm_12_3_1);
  assign argmax_else_acc_nl = nl_argmax_else_acc_nl[10:0];
  assign argmax_else_if_argmax_else_if_argmax_else_if_nor_nl = ~((readslicef_11_1_10(argmax_else_aif_acc_nl))
      | (readslicef_11_1_10(argmax_else_acc_nl)));
  assign argmax_else_mux_nl = MUX_v_2_2_2(2'b01, 2'b10, argmax_else_if_argmax_else_if_argmax_else_if_nor_nl);
  assign nl_argmax_aif_acc_nl = conv_s2u_10_11(Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_itm_12_3_1)
      - conv_s2u_10_11(Accum1_1_58_Accum2_1_3_Accum2_1_acc_1_itm_12_3_1);
  assign argmax_aif_acc_nl = nl_argmax_aif_acc_nl[10:0];
  assign nl_argmax_acc_nl = conv_s2u_10_11(Accum1_1_58_Accum2_1_1_Accum2_1_acc_1_itm_12_3_1)
      - conv_s2u_10_11(Accum1_1_58_Accum2_1_2_Accum2_1_acc_1_itm_12_3_1);
  assign argmax_acc_nl = nl_argmax_acc_nl[10:0];
  assign argmax_if_argmax_if_argmax_if_nor_nl = ~((readslicef_11_1_10(argmax_aif_acc_nl))
      | (readslicef_11_1_10(argmax_acc_nl)));

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] readslicef_13_10_3;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_13_10_3 = tmp[9:0];
  end
  endfunction


  function automatic [8:0] readslicef_15_9_6;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_15_9_6 = tmp[8:0];
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_5_9 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_9 = {{4{vector[4]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_9_13 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_13 = {{4{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_10_13 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_13 = {{3{vector[9]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    myproject
// ------------------------------------------------------------------


module myproject (
  clk, rst, input_1_rsc_dat, layer7_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [95:0] input_1_rsc_dat;
  output [1:0] layer7_out_rsc_dat;
  input [4639:0] w2_rsc_dat;
  input [289:0] b2_rsc_dat;
  input [869:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  converterBlock_myproject_core myproject_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .w2_rsc_dat(w2_rsc_dat),
      .b2_rsc_dat(b2_rsc_dat),
      .w5_rsc_dat(w5_rsc_dat),
      .b5_rsc_dat(b5_rsc_dat)
    );
endmodule



