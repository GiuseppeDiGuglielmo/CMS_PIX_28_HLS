
//------> ./myproject_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module converterBlock_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./myproject_ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module converterBlock_ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> ./myproject.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2022.1_1/994485 Production Release
//  HLS Date:       Mon May  9 08:51:12 PDT 2022
// 
//  Generated by:   giuseppe@ml4asic01
//  Generated date: Tue Dec 13 20:57:48 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    converterBlock_myproject_core
// ------------------------------------------------------------------


module converterBlock_myproject_core (
  clk, rst, input_1_rsc_dat, layer7_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [95:0] input_1_rsc_dat;
  output [1:0] layer7_out_rsc_dat;
  input [5119:0] w2_rsc_dat;
  input [319:0] b2_rsc_dat;
  input [959:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;


  // Interconnect Declarations
  wire [95:0] input_1_rsci_idat;
  reg [1:0] layer7_out_rsci_idat;
  wire [5119:0] w2_rsci_idat;
  wire [319:0] b2_rsci_idat;
  wire [959:0] w5_rsci_idat;
  wire [14:0] b5_rsci_idat;
  wire [15:0] Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1;
  wire [21:0] nl_Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1;
  wire [11:0] Accum2_acc_127_psp_sva_1;
  wire [12:0] nl_Accum2_acc_127_psp_sva_1;
  wire [11:0] Accum2_acc_126_psp_sva_1;
  wire [12:0] nl_Accum2_acc_126_psp_sva_1;
  wire [11:0] Accum2_acc_125_psp_sva_1;
  wire [12:0] nl_Accum2_acc_125_psp_sva_1;
  wire [11:0] Accum2_acc_124_psp_sva_1;
  wire [12:0] nl_Accum2_acc_124_psp_sva_1;
  wire [11:0] Accum2_acc_123_psp_sva_1;
  wire [12:0] nl_Accum2_acc_123_psp_sva_1;
  wire [11:0] Accum2_acc_122_psp_sva_1;
  wire [12:0] nl_Accum2_acc_122_psp_sva_1;
  wire [11:0] Accum2_acc_121_psp_sva_1;
  wire [12:0] nl_Accum2_acc_121_psp_sva_1;
  wire [11:0] Accum2_acc_120_psp_sva_1;
  wire [12:0] nl_Accum2_acc_120_psp_sva_1;
  wire [11:0] Accum2_acc_119_psp_sva_1;
  wire [12:0] nl_Accum2_acc_119_psp_sva_1;
  wire [11:0] Accum2_acc_118_psp_sva_1;
  wire [12:0] nl_Accum2_acc_118_psp_sva_1;
  wire [11:0] Accum2_acc_117_psp_sva_1;
  wire [12:0] nl_Accum2_acc_117_psp_sva_1;
  wire [11:0] Accum2_acc_116_psp_sva_1;
  wire [12:0] nl_Accum2_acc_116_psp_sva_1;
  wire [11:0] Accum2_acc_115_psp_sva_1;
  wire [12:0] nl_Accum2_acc_115_psp_sva_1;
  wire [11:0] Accum2_acc_114_psp_sva_1;
  wire [12:0] nl_Accum2_acc_114_psp_sva_1;
  wire [11:0] Accum2_acc_113_psp_sva_1;
  wire [12:0] nl_Accum2_acc_113_psp_sva_1;
  wire [11:0] Accum2_acc_112_psp_sva_1;
  wire [12:0] nl_Accum2_acc_112_psp_sva_1;
  wire [11:0] Accum2_acc_111_psp_sva_1;
  wire [12:0] nl_Accum2_acc_111_psp_sva_1;
  wire [11:0] Accum2_acc_110_psp_sva_1;
  wire [12:0] nl_Accum2_acc_110_psp_sva_1;
  wire [11:0] Accum2_acc_109_psp_sva_1;
  wire [12:0] nl_Accum2_acc_109_psp_sva_1;
  wire [11:0] Accum2_acc_108_psp_sva_1;
  wire [12:0] nl_Accum2_acc_108_psp_sva_1;
  wire [11:0] Accum2_acc_107_psp_sva_1;
  wire [12:0] nl_Accum2_acc_107_psp_sva_1;
  wire [11:0] Accum2_acc_106_psp_sva_1;
  wire [12:0] nl_Accum2_acc_106_psp_sva_1;
  wire [11:0] Accum2_acc_105_psp_sva_1;
  wire [12:0] nl_Accum2_acc_105_psp_sva_1;
  wire [11:0] Accum2_acc_104_psp_sva_1;
  wire [12:0] nl_Accum2_acc_104_psp_sva_1;
  wire [11:0] Accum2_acc_103_psp_sva_1;
  wire [12:0] nl_Accum2_acc_103_psp_sva_1;
  wire [11:0] Accum2_acc_102_psp_sva_1;
  wire [12:0] nl_Accum2_acc_102_psp_sva_1;
  wire [11:0] Accum2_acc_101_psp_sva_1;
  wire [12:0] nl_Accum2_acc_101_psp_sva_1;
  wire [11:0] Accum2_acc_100_psp_sva_1;
  wire [12:0] nl_Accum2_acc_100_psp_sva_1;
  wire [11:0] Accum2_acc_99_psp_sva_1;
  wire [12:0] nl_Accum2_acc_99_psp_sva_1;
  wire [11:0] Accum2_acc_98_psp_sva_1;
  wire [12:0] nl_Accum2_acc_98_psp_sva_1;
  wire [11:0] Accum2_acc_97_psp_sva_1;
  wire [12:0] nl_Accum2_acc_97_psp_sva_1;
  wire [11:0] Accum2_acc_96_psp_sva_1;
  wire [12:0] nl_Accum2_acc_96_psp_sva_1;
  wire [11:0] Accum2_acc_95_psp_sva_1;
  wire [12:0] nl_Accum2_acc_95_psp_sva_1;
  wire [11:0] Accum2_acc_94_psp_sva_1;
  wire [12:0] nl_Accum2_acc_94_psp_sva_1;
  wire [11:0] Accum2_acc_93_psp_sva_1;
  wire [12:0] nl_Accum2_acc_93_psp_sva_1;
  wire [11:0] Accum2_acc_92_psp_sva_1;
  wire [12:0] nl_Accum2_acc_92_psp_sva_1;
  wire [11:0] Accum2_acc_91_psp_sva_1;
  wire [12:0] nl_Accum2_acc_91_psp_sva_1;
  wire [11:0] Accum2_acc_90_psp_sva_1;
  wire [12:0] nl_Accum2_acc_90_psp_sva_1;
  wire [11:0] Accum2_acc_89_psp_sva_1;
  wire [12:0] nl_Accum2_acc_89_psp_sva_1;
  wire [11:0] Accum2_acc_88_psp_sva_1;
  wire [12:0] nl_Accum2_acc_88_psp_sva_1;
  wire [11:0] Accum2_acc_87_psp_sva_1;
  wire [12:0] nl_Accum2_acc_87_psp_sva_1;
  wire [11:0] Accum2_acc_86_psp_sva_1;
  wire [12:0] nl_Accum2_acc_86_psp_sva_1;
  wire [11:0] Accum2_acc_85_psp_sva_1;
  wire [12:0] nl_Accum2_acc_85_psp_sva_1;
  wire [11:0] Accum2_acc_84_psp_sva_1;
  wire [12:0] nl_Accum2_acc_84_psp_sva_1;
  wire [11:0] Accum2_acc_83_psp_sva_1;
  wire [12:0] nl_Accum2_acc_83_psp_sva_1;
  wire [11:0] Accum2_acc_82_psp_sva_1;
  wire [12:0] nl_Accum2_acc_82_psp_sva_1;
  wire [11:0] Accum2_acc_81_psp_sva_1;
  wire [12:0] nl_Accum2_acc_81_psp_sva_1;
  wire [11:0] Accum2_acc_80_psp_sva_1;
  wire [12:0] nl_Accum2_acc_80_psp_sva_1;
  wire [11:0] Accum2_acc_79_psp_sva_1;
  wire [12:0] nl_Accum2_acc_79_psp_sva_1;
  wire [11:0] Accum2_acc_78_psp_sva_1;
  wire [12:0] nl_Accum2_acc_78_psp_sva_1;
  wire [11:0] Accum2_acc_77_psp_sva_1;
  wire [12:0] nl_Accum2_acc_77_psp_sva_1;
  wire [11:0] Accum2_acc_76_psp_sva_1;
  wire [12:0] nl_Accum2_acc_76_psp_sva_1;
  wire [11:0] Accum2_acc_75_psp_sva_1;
  wire [12:0] nl_Accum2_acc_75_psp_sva_1;
  wire [11:0] Accum2_acc_74_psp_sva_1;
  wire [12:0] nl_Accum2_acc_74_psp_sva_1;
  wire [11:0] Accum2_acc_73_psp_sva_1;
  wire [12:0] nl_Accum2_acc_73_psp_sva_1;
  wire [11:0] Accum2_acc_72_psp_sva_1;
  wire [12:0] nl_Accum2_acc_72_psp_sva_1;
  wire [11:0] Accum2_acc_71_psp_sva_1;
  wire [12:0] nl_Accum2_acc_71_psp_sva_1;
  wire [11:0] Accum2_acc_70_psp_sva_1;
  wire [12:0] nl_Accum2_acc_70_psp_sva_1;
  wire [11:0] Accum2_acc_69_psp_sva_1;
  wire [12:0] nl_Accum2_acc_69_psp_sva_1;
  wire [11:0] Accum2_acc_68_psp_sva_1;
  wire [12:0] nl_Accum2_acc_68_psp_sva_1;
  wire [11:0] Accum2_acc_67_psp_sva_1;
  wire [12:0] nl_Accum2_acc_67_psp_sva_1;
  wire [11:0] Accum2_acc_66_psp_sva_1;
  wire [12:0] nl_Accum2_acc_66_psp_sva_1;
  wire [11:0] Accum2_acc_65_psp_sva_1;
  wire [12:0] nl_Accum2_acc_65_psp_sva_1;
  wire [15:0] Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1;
  wire [21:0] nl_Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1;
  wire [15:0] Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1;
  wire [21:0] nl_Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1;
  wire [11:0] layer3_out_0_15_4_sva_1;
  wire [12:0] nl_layer3_out_0_15_4_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire layer4_out_0_2_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_8_6;
  wire layer4_out_conc_4_9;
  wire [2:0] layer4_out_conc_4_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_6;
  wire nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9;
  wire [2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_6;
  wire [8:0] Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1;
  wire [8:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1;
  wire [8:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_12_1;
  wire operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_12_1;

  wire[1:0] argmax_else_mux_nl;
  wire argmax_else_if_argmax_else_if_argmax_else_if_nor_nl;
  wire[15:0] argmax_else_aif_acc_nl;
  wire[16:0] nl_argmax_else_aif_acc_nl;
  wire[15:0] argmax_else_acc_nl;
  wire[16:0] nl_argmax_else_acc_nl;
  wire argmax_if_argmax_if_argmax_if_nor_nl;
  wire[15:0] argmax_aif_acc_nl;
  wire[16:0] nl_argmax_aif_acc_nl;
  wire[15:0] argmax_acc_nl;
  wire[16:0] nl_argmax_acc_nl;
  wire[11:0] Accum2_acc_1968_nl;
  wire[14:0] nl_Accum2_acc_1968_nl;
  wire[11:0] Accum2_acc_1965_nl;
  wire[13:0] nl_Accum2_acc_1965_nl;
  wire[10:0] Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1954_nl;
  wire[11:0] nl_Accum2_acc_1954_nl;
  wire[10:0] Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1967_nl;
  wire[14:0] nl_Accum2_acc_1967_nl;
  wire[11:0] Accum2_acc_1963_nl;
  wire[13:0] nl_Accum2_acc_1963_nl;
  wire[10:0] Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_nl;
  wire[14:0] nl_Accum2_acc_nl;
  wire[11:0] Accum2_acc_1020_nl;
  wire[13:0] nl_Accum2_acc_1020_nl;
  wire[10:0] Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1017_nl;
  wire[11:0] nl_Accum2_acc_1017_nl;
  wire[10:0] Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1022_nl;
  wire[14:0] nl_Accum2_acc_1022_nl;
  wire[11:0] Accum2_acc_1018_nl;
  wire[13:0] nl_Accum2_acc_1018_nl;
  wire[10:0] Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1038_nl;
  wire[14:0] nl_Accum2_acc_1038_nl;
  wire[11:0] Accum2_acc_1035_nl;
  wire[13:0] nl_Accum2_acc_1035_nl;
  wire[10:0] Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1024_nl;
  wire[11:0] nl_Accum2_acc_1024_nl;
  wire[10:0] Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1037_nl;
  wire[14:0] nl_Accum2_acc_1037_nl;
  wire[11:0] Accum2_acc_1033_nl;
  wire[13:0] nl_Accum2_acc_1033_nl;
  wire[10:0] Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1053_nl;
  wire[14:0] nl_Accum2_acc_1053_nl;
  wire[11:0] Accum2_acc_1050_nl;
  wire[13:0] nl_Accum2_acc_1050_nl;
  wire[10:0] Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1039_nl;
  wire[11:0] nl_Accum2_acc_1039_nl;
  wire[10:0] Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1052_nl;
  wire[14:0] nl_Accum2_acc_1052_nl;
  wire[11:0] Accum2_acc_1048_nl;
  wire[13:0] nl_Accum2_acc_1048_nl;
  wire[10:0] Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1068_nl;
  wire[14:0] nl_Accum2_acc_1068_nl;
  wire[11:0] Accum2_acc_1065_nl;
  wire[13:0] nl_Accum2_acc_1065_nl;
  wire[10:0] Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1054_nl;
  wire[11:0] nl_Accum2_acc_1054_nl;
  wire[10:0] Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1067_nl;
  wire[14:0] nl_Accum2_acc_1067_nl;
  wire[11:0] Accum2_acc_1063_nl;
  wire[13:0] nl_Accum2_acc_1063_nl;
  wire[10:0] Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1083_nl;
  wire[14:0] nl_Accum2_acc_1083_nl;
  wire[11:0] Accum2_acc_1080_nl;
  wire[13:0] nl_Accum2_acc_1080_nl;
  wire[10:0] Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1069_nl;
  wire[11:0] nl_Accum2_acc_1069_nl;
  wire[10:0] Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1082_nl;
  wire[14:0] nl_Accum2_acc_1082_nl;
  wire[11:0] Accum2_acc_1078_nl;
  wire[13:0] nl_Accum2_acc_1078_nl;
  wire[10:0] Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1098_nl;
  wire[14:0] nl_Accum2_acc_1098_nl;
  wire[11:0] Accum2_acc_1095_nl;
  wire[13:0] nl_Accum2_acc_1095_nl;
  wire[10:0] Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1084_nl;
  wire[11:0] nl_Accum2_acc_1084_nl;
  wire[10:0] Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1097_nl;
  wire[14:0] nl_Accum2_acc_1097_nl;
  wire[11:0] Accum2_acc_1093_nl;
  wire[13:0] nl_Accum2_acc_1093_nl;
  wire[10:0] Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1113_nl;
  wire[14:0] nl_Accum2_acc_1113_nl;
  wire[11:0] Accum2_acc_1110_nl;
  wire[13:0] nl_Accum2_acc_1110_nl;
  wire[10:0] Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1099_nl;
  wire[11:0] nl_Accum2_acc_1099_nl;
  wire[10:0] Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1112_nl;
  wire[14:0] nl_Accum2_acc_1112_nl;
  wire[11:0] Accum2_acc_1108_nl;
  wire[13:0] nl_Accum2_acc_1108_nl;
  wire[10:0] Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1128_nl;
  wire[14:0] nl_Accum2_acc_1128_nl;
  wire[11:0] Accum2_acc_1125_nl;
  wire[13:0] nl_Accum2_acc_1125_nl;
  wire[10:0] Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1114_nl;
  wire[11:0] nl_Accum2_acc_1114_nl;
  wire[10:0] Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1127_nl;
  wire[14:0] nl_Accum2_acc_1127_nl;
  wire[11:0] Accum2_acc_1123_nl;
  wire[13:0] nl_Accum2_acc_1123_nl;
  wire[10:0] Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1143_nl;
  wire[14:0] nl_Accum2_acc_1143_nl;
  wire[11:0] Accum2_acc_1140_nl;
  wire[13:0] nl_Accum2_acc_1140_nl;
  wire[10:0] Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1129_nl;
  wire[11:0] nl_Accum2_acc_1129_nl;
  wire[10:0] Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1142_nl;
  wire[14:0] nl_Accum2_acc_1142_nl;
  wire[11:0] Accum2_acc_1138_nl;
  wire[13:0] nl_Accum2_acc_1138_nl;
  wire[10:0] Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1158_nl;
  wire[14:0] nl_Accum2_acc_1158_nl;
  wire[11:0] Accum2_acc_1155_nl;
  wire[13:0] nl_Accum2_acc_1155_nl;
  wire[10:0] Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1144_nl;
  wire[11:0] nl_Accum2_acc_1144_nl;
  wire[10:0] Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1157_nl;
  wire[14:0] nl_Accum2_acc_1157_nl;
  wire[11:0] Accum2_acc_1153_nl;
  wire[13:0] nl_Accum2_acc_1153_nl;
  wire[10:0] Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1173_nl;
  wire[14:0] nl_Accum2_acc_1173_nl;
  wire[11:0] Accum2_acc_1170_nl;
  wire[13:0] nl_Accum2_acc_1170_nl;
  wire[10:0] Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1159_nl;
  wire[11:0] nl_Accum2_acc_1159_nl;
  wire[10:0] Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1172_nl;
  wire[14:0] nl_Accum2_acc_1172_nl;
  wire[11:0] Accum2_acc_1168_nl;
  wire[13:0] nl_Accum2_acc_1168_nl;
  wire[10:0] Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1188_nl;
  wire[14:0] nl_Accum2_acc_1188_nl;
  wire[11:0] Accum2_acc_1185_nl;
  wire[13:0] nl_Accum2_acc_1185_nl;
  wire[10:0] Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1174_nl;
  wire[11:0] nl_Accum2_acc_1174_nl;
  wire[10:0] Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1187_nl;
  wire[14:0] nl_Accum2_acc_1187_nl;
  wire[11:0] Accum2_acc_1183_nl;
  wire[13:0] nl_Accum2_acc_1183_nl;
  wire[10:0] Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1203_nl;
  wire[14:0] nl_Accum2_acc_1203_nl;
  wire[11:0] Accum2_acc_1200_nl;
  wire[13:0] nl_Accum2_acc_1200_nl;
  wire[10:0] Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1189_nl;
  wire[11:0] nl_Accum2_acc_1189_nl;
  wire[10:0] Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1202_nl;
  wire[14:0] nl_Accum2_acc_1202_nl;
  wire[11:0] Accum2_acc_1198_nl;
  wire[13:0] nl_Accum2_acc_1198_nl;
  wire[10:0] Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1218_nl;
  wire[14:0] nl_Accum2_acc_1218_nl;
  wire[11:0] Accum2_acc_1215_nl;
  wire[13:0] nl_Accum2_acc_1215_nl;
  wire[10:0] Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1204_nl;
  wire[11:0] nl_Accum2_acc_1204_nl;
  wire[10:0] Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1217_nl;
  wire[14:0] nl_Accum2_acc_1217_nl;
  wire[11:0] Accum2_acc_1213_nl;
  wire[13:0] nl_Accum2_acc_1213_nl;
  wire[10:0] Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1233_nl;
  wire[14:0] nl_Accum2_acc_1233_nl;
  wire[11:0] Accum2_acc_1230_nl;
  wire[13:0] nl_Accum2_acc_1230_nl;
  wire[10:0] Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1219_nl;
  wire[11:0] nl_Accum2_acc_1219_nl;
  wire[10:0] Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1232_nl;
  wire[14:0] nl_Accum2_acc_1232_nl;
  wire[11:0] Accum2_acc_1228_nl;
  wire[13:0] nl_Accum2_acc_1228_nl;
  wire[10:0] Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1248_nl;
  wire[14:0] nl_Accum2_acc_1248_nl;
  wire[11:0] Accum2_acc_1245_nl;
  wire[13:0] nl_Accum2_acc_1245_nl;
  wire[10:0] Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1234_nl;
  wire[11:0] nl_Accum2_acc_1234_nl;
  wire[10:0] Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1247_nl;
  wire[14:0] nl_Accum2_acc_1247_nl;
  wire[11:0] Accum2_acc_1243_nl;
  wire[13:0] nl_Accum2_acc_1243_nl;
  wire[10:0] Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1263_nl;
  wire[14:0] nl_Accum2_acc_1263_nl;
  wire[11:0] Accum2_acc_1260_nl;
  wire[13:0] nl_Accum2_acc_1260_nl;
  wire[10:0] Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1249_nl;
  wire[11:0] nl_Accum2_acc_1249_nl;
  wire[10:0] Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1262_nl;
  wire[14:0] nl_Accum2_acc_1262_nl;
  wire[11:0] Accum2_acc_1258_nl;
  wire[13:0] nl_Accum2_acc_1258_nl;
  wire[10:0] Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1278_nl;
  wire[14:0] nl_Accum2_acc_1278_nl;
  wire[11:0] Accum2_acc_1275_nl;
  wire[13:0] nl_Accum2_acc_1275_nl;
  wire[10:0] Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1264_nl;
  wire[11:0] nl_Accum2_acc_1264_nl;
  wire[10:0] Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1277_nl;
  wire[14:0] nl_Accum2_acc_1277_nl;
  wire[11:0] Accum2_acc_1273_nl;
  wire[13:0] nl_Accum2_acc_1273_nl;
  wire[10:0] Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1293_nl;
  wire[14:0] nl_Accum2_acc_1293_nl;
  wire[11:0] Accum2_acc_1290_nl;
  wire[13:0] nl_Accum2_acc_1290_nl;
  wire[10:0] Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1279_nl;
  wire[11:0] nl_Accum2_acc_1279_nl;
  wire[10:0] Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1292_nl;
  wire[14:0] nl_Accum2_acc_1292_nl;
  wire[11:0] Accum2_acc_1288_nl;
  wire[13:0] nl_Accum2_acc_1288_nl;
  wire[10:0] Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1308_nl;
  wire[14:0] nl_Accum2_acc_1308_nl;
  wire[11:0] Accum2_acc_1305_nl;
  wire[13:0] nl_Accum2_acc_1305_nl;
  wire[10:0] Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1294_nl;
  wire[11:0] nl_Accum2_acc_1294_nl;
  wire[10:0] Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1307_nl;
  wire[14:0] nl_Accum2_acc_1307_nl;
  wire[11:0] Accum2_acc_1303_nl;
  wire[13:0] nl_Accum2_acc_1303_nl;
  wire[10:0] Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1323_nl;
  wire[14:0] nl_Accum2_acc_1323_nl;
  wire[11:0] Accum2_acc_1320_nl;
  wire[13:0] nl_Accum2_acc_1320_nl;
  wire[10:0] Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1309_nl;
  wire[11:0] nl_Accum2_acc_1309_nl;
  wire[10:0] Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1322_nl;
  wire[14:0] nl_Accum2_acc_1322_nl;
  wire[11:0] Accum2_acc_1318_nl;
  wire[13:0] nl_Accum2_acc_1318_nl;
  wire[10:0] Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1338_nl;
  wire[14:0] nl_Accum2_acc_1338_nl;
  wire[11:0] Accum2_acc_1335_nl;
  wire[13:0] nl_Accum2_acc_1335_nl;
  wire[10:0] Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1324_nl;
  wire[11:0] nl_Accum2_acc_1324_nl;
  wire[10:0] Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1337_nl;
  wire[14:0] nl_Accum2_acc_1337_nl;
  wire[11:0] Accum2_acc_1333_nl;
  wire[13:0] nl_Accum2_acc_1333_nl;
  wire[10:0] Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1353_nl;
  wire[14:0] nl_Accum2_acc_1353_nl;
  wire[11:0] Accum2_acc_1350_nl;
  wire[13:0] nl_Accum2_acc_1350_nl;
  wire[10:0] Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1339_nl;
  wire[11:0] nl_Accum2_acc_1339_nl;
  wire[10:0] Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1352_nl;
  wire[14:0] nl_Accum2_acc_1352_nl;
  wire[11:0] Accum2_acc_1348_nl;
  wire[13:0] nl_Accum2_acc_1348_nl;
  wire[10:0] Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1368_nl;
  wire[14:0] nl_Accum2_acc_1368_nl;
  wire[11:0] Accum2_acc_1365_nl;
  wire[13:0] nl_Accum2_acc_1365_nl;
  wire[10:0] Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1354_nl;
  wire[11:0] nl_Accum2_acc_1354_nl;
  wire[10:0] Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1367_nl;
  wire[14:0] nl_Accum2_acc_1367_nl;
  wire[11:0] Accum2_acc_1363_nl;
  wire[13:0] nl_Accum2_acc_1363_nl;
  wire[10:0] Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1383_nl;
  wire[14:0] nl_Accum2_acc_1383_nl;
  wire[11:0] Accum2_acc_1380_nl;
  wire[13:0] nl_Accum2_acc_1380_nl;
  wire[10:0] Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1369_nl;
  wire[11:0] nl_Accum2_acc_1369_nl;
  wire[10:0] Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1382_nl;
  wire[14:0] nl_Accum2_acc_1382_nl;
  wire[11:0] Accum2_acc_1378_nl;
  wire[13:0] nl_Accum2_acc_1378_nl;
  wire[10:0] Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1398_nl;
  wire[14:0] nl_Accum2_acc_1398_nl;
  wire[11:0] Accum2_acc_1395_nl;
  wire[13:0] nl_Accum2_acc_1395_nl;
  wire[10:0] Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1384_nl;
  wire[11:0] nl_Accum2_acc_1384_nl;
  wire[10:0] Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1397_nl;
  wire[14:0] nl_Accum2_acc_1397_nl;
  wire[11:0] Accum2_acc_1393_nl;
  wire[13:0] nl_Accum2_acc_1393_nl;
  wire[10:0] Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1413_nl;
  wire[14:0] nl_Accum2_acc_1413_nl;
  wire[11:0] Accum2_acc_1410_nl;
  wire[13:0] nl_Accum2_acc_1410_nl;
  wire[10:0] Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1399_nl;
  wire[11:0] nl_Accum2_acc_1399_nl;
  wire[10:0] Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1412_nl;
  wire[14:0] nl_Accum2_acc_1412_nl;
  wire[11:0] Accum2_acc_1408_nl;
  wire[13:0] nl_Accum2_acc_1408_nl;
  wire[10:0] Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1428_nl;
  wire[14:0] nl_Accum2_acc_1428_nl;
  wire[11:0] Accum2_acc_1425_nl;
  wire[13:0] nl_Accum2_acc_1425_nl;
  wire[10:0] Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1414_nl;
  wire[11:0] nl_Accum2_acc_1414_nl;
  wire[10:0] Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1427_nl;
  wire[14:0] nl_Accum2_acc_1427_nl;
  wire[11:0] Accum2_acc_1423_nl;
  wire[13:0] nl_Accum2_acc_1423_nl;
  wire[10:0] Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1443_nl;
  wire[14:0] nl_Accum2_acc_1443_nl;
  wire[11:0] Accum2_acc_1440_nl;
  wire[13:0] nl_Accum2_acc_1440_nl;
  wire[10:0] Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1429_nl;
  wire[11:0] nl_Accum2_acc_1429_nl;
  wire[10:0] Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1442_nl;
  wire[14:0] nl_Accum2_acc_1442_nl;
  wire[11:0] Accum2_acc_1438_nl;
  wire[13:0] nl_Accum2_acc_1438_nl;
  wire[10:0] Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1458_nl;
  wire[14:0] nl_Accum2_acc_1458_nl;
  wire[11:0] Accum2_acc_1455_nl;
  wire[13:0] nl_Accum2_acc_1455_nl;
  wire[10:0] Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1444_nl;
  wire[11:0] nl_Accum2_acc_1444_nl;
  wire[10:0] Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1457_nl;
  wire[14:0] nl_Accum2_acc_1457_nl;
  wire[11:0] Accum2_acc_1453_nl;
  wire[13:0] nl_Accum2_acc_1453_nl;
  wire[10:0] Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1473_nl;
  wire[14:0] nl_Accum2_acc_1473_nl;
  wire[11:0] Accum2_acc_1470_nl;
  wire[13:0] nl_Accum2_acc_1470_nl;
  wire[10:0] Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1459_nl;
  wire[11:0] nl_Accum2_acc_1459_nl;
  wire[10:0] Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1472_nl;
  wire[14:0] nl_Accum2_acc_1472_nl;
  wire[11:0] Accum2_acc_1468_nl;
  wire[13:0] nl_Accum2_acc_1468_nl;
  wire[10:0] Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1488_nl;
  wire[14:0] nl_Accum2_acc_1488_nl;
  wire[11:0] Accum2_acc_1485_nl;
  wire[13:0] nl_Accum2_acc_1485_nl;
  wire[10:0] Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1474_nl;
  wire[11:0] nl_Accum2_acc_1474_nl;
  wire[10:0] Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1487_nl;
  wire[14:0] nl_Accum2_acc_1487_nl;
  wire[11:0] Accum2_acc_1483_nl;
  wire[13:0] nl_Accum2_acc_1483_nl;
  wire[10:0] Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1503_nl;
  wire[14:0] nl_Accum2_acc_1503_nl;
  wire[11:0] Accum2_acc_1500_nl;
  wire[13:0] nl_Accum2_acc_1500_nl;
  wire[10:0] Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1489_nl;
  wire[11:0] nl_Accum2_acc_1489_nl;
  wire[10:0] Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1502_nl;
  wire[14:0] nl_Accum2_acc_1502_nl;
  wire[11:0] Accum2_acc_1498_nl;
  wire[13:0] nl_Accum2_acc_1498_nl;
  wire[10:0] Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1518_nl;
  wire[14:0] nl_Accum2_acc_1518_nl;
  wire[11:0] Accum2_acc_1515_nl;
  wire[13:0] nl_Accum2_acc_1515_nl;
  wire[10:0] Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1504_nl;
  wire[11:0] nl_Accum2_acc_1504_nl;
  wire[10:0] Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1517_nl;
  wire[14:0] nl_Accum2_acc_1517_nl;
  wire[11:0] Accum2_acc_1513_nl;
  wire[13:0] nl_Accum2_acc_1513_nl;
  wire[10:0] Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1533_nl;
  wire[14:0] nl_Accum2_acc_1533_nl;
  wire[11:0] Accum2_acc_1530_nl;
  wire[13:0] nl_Accum2_acc_1530_nl;
  wire[10:0] Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1519_nl;
  wire[11:0] nl_Accum2_acc_1519_nl;
  wire[10:0] Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1532_nl;
  wire[14:0] nl_Accum2_acc_1532_nl;
  wire[11:0] Accum2_acc_1528_nl;
  wire[13:0] nl_Accum2_acc_1528_nl;
  wire[10:0] Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1548_nl;
  wire[14:0] nl_Accum2_acc_1548_nl;
  wire[11:0] Accum2_acc_1545_nl;
  wire[13:0] nl_Accum2_acc_1545_nl;
  wire[10:0] Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1534_nl;
  wire[11:0] nl_Accum2_acc_1534_nl;
  wire[10:0] Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1547_nl;
  wire[14:0] nl_Accum2_acc_1547_nl;
  wire[11:0] Accum2_acc_1543_nl;
  wire[13:0] nl_Accum2_acc_1543_nl;
  wire[10:0] Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1563_nl;
  wire[14:0] nl_Accum2_acc_1563_nl;
  wire[11:0] Accum2_acc_1560_nl;
  wire[13:0] nl_Accum2_acc_1560_nl;
  wire[10:0] Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1549_nl;
  wire[11:0] nl_Accum2_acc_1549_nl;
  wire[10:0] Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1562_nl;
  wire[14:0] nl_Accum2_acc_1562_nl;
  wire[11:0] Accum2_acc_1558_nl;
  wire[13:0] nl_Accum2_acc_1558_nl;
  wire[10:0] Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1578_nl;
  wire[14:0] nl_Accum2_acc_1578_nl;
  wire[11:0] Accum2_acc_1575_nl;
  wire[13:0] nl_Accum2_acc_1575_nl;
  wire[10:0] Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1564_nl;
  wire[11:0] nl_Accum2_acc_1564_nl;
  wire[10:0] Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1577_nl;
  wire[14:0] nl_Accum2_acc_1577_nl;
  wire[11:0] Accum2_acc_1573_nl;
  wire[13:0] nl_Accum2_acc_1573_nl;
  wire[10:0] Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1593_nl;
  wire[14:0] nl_Accum2_acc_1593_nl;
  wire[11:0] Accum2_acc_1590_nl;
  wire[13:0] nl_Accum2_acc_1590_nl;
  wire[10:0] Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1579_nl;
  wire[11:0] nl_Accum2_acc_1579_nl;
  wire[10:0] Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1592_nl;
  wire[14:0] nl_Accum2_acc_1592_nl;
  wire[11:0] Accum2_acc_1588_nl;
  wire[13:0] nl_Accum2_acc_1588_nl;
  wire[10:0] Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1608_nl;
  wire[14:0] nl_Accum2_acc_1608_nl;
  wire[11:0] Accum2_acc_1605_nl;
  wire[13:0] nl_Accum2_acc_1605_nl;
  wire[10:0] Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1594_nl;
  wire[11:0] nl_Accum2_acc_1594_nl;
  wire[10:0] Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1607_nl;
  wire[14:0] nl_Accum2_acc_1607_nl;
  wire[11:0] Accum2_acc_1603_nl;
  wire[13:0] nl_Accum2_acc_1603_nl;
  wire[10:0] Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1623_nl;
  wire[14:0] nl_Accum2_acc_1623_nl;
  wire[11:0] Accum2_acc_1620_nl;
  wire[13:0] nl_Accum2_acc_1620_nl;
  wire[10:0] Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1609_nl;
  wire[11:0] nl_Accum2_acc_1609_nl;
  wire[10:0] Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1622_nl;
  wire[14:0] nl_Accum2_acc_1622_nl;
  wire[11:0] Accum2_acc_1618_nl;
  wire[13:0] nl_Accum2_acc_1618_nl;
  wire[10:0] Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1638_nl;
  wire[14:0] nl_Accum2_acc_1638_nl;
  wire[11:0] Accum2_acc_1635_nl;
  wire[13:0] nl_Accum2_acc_1635_nl;
  wire[10:0] Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1624_nl;
  wire[11:0] nl_Accum2_acc_1624_nl;
  wire[10:0] Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1637_nl;
  wire[14:0] nl_Accum2_acc_1637_nl;
  wire[11:0] Accum2_acc_1633_nl;
  wire[13:0] nl_Accum2_acc_1633_nl;
  wire[10:0] Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1653_nl;
  wire[14:0] nl_Accum2_acc_1653_nl;
  wire[11:0] Accum2_acc_1650_nl;
  wire[13:0] nl_Accum2_acc_1650_nl;
  wire[10:0] Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1639_nl;
  wire[11:0] nl_Accum2_acc_1639_nl;
  wire[10:0] Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1652_nl;
  wire[14:0] nl_Accum2_acc_1652_nl;
  wire[11:0] Accum2_acc_1648_nl;
  wire[13:0] nl_Accum2_acc_1648_nl;
  wire[10:0] Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1668_nl;
  wire[14:0] nl_Accum2_acc_1668_nl;
  wire[11:0] Accum2_acc_1665_nl;
  wire[13:0] nl_Accum2_acc_1665_nl;
  wire[10:0] Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1654_nl;
  wire[11:0] nl_Accum2_acc_1654_nl;
  wire[10:0] Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1667_nl;
  wire[14:0] nl_Accum2_acc_1667_nl;
  wire[11:0] Accum2_acc_1663_nl;
  wire[13:0] nl_Accum2_acc_1663_nl;
  wire[10:0] Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1683_nl;
  wire[14:0] nl_Accum2_acc_1683_nl;
  wire[11:0] Accum2_acc_1680_nl;
  wire[13:0] nl_Accum2_acc_1680_nl;
  wire[10:0] Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1669_nl;
  wire[11:0] nl_Accum2_acc_1669_nl;
  wire[10:0] Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1682_nl;
  wire[14:0] nl_Accum2_acc_1682_nl;
  wire[11:0] Accum2_acc_1678_nl;
  wire[13:0] nl_Accum2_acc_1678_nl;
  wire[10:0] Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1698_nl;
  wire[14:0] nl_Accum2_acc_1698_nl;
  wire[11:0] Accum2_acc_1695_nl;
  wire[13:0] nl_Accum2_acc_1695_nl;
  wire[10:0] Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1684_nl;
  wire[11:0] nl_Accum2_acc_1684_nl;
  wire[10:0] Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1697_nl;
  wire[14:0] nl_Accum2_acc_1697_nl;
  wire[11:0] Accum2_acc_1693_nl;
  wire[13:0] nl_Accum2_acc_1693_nl;
  wire[10:0] Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1713_nl;
  wire[14:0] nl_Accum2_acc_1713_nl;
  wire[11:0] Accum2_acc_1710_nl;
  wire[13:0] nl_Accum2_acc_1710_nl;
  wire[10:0] Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1699_nl;
  wire[11:0] nl_Accum2_acc_1699_nl;
  wire[10:0] Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1712_nl;
  wire[14:0] nl_Accum2_acc_1712_nl;
  wire[11:0] Accum2_acc_1708_nl;
  wire[13:0] nl_Accum2_acc_1708_nl;
  wire[10:0] Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1728_nl;
  wire[14:0] nl_Accum2_acc_1728_nl;
  wire[11:0] Accum2_acc_1725_nl;
  wire[13:0] nl_Accum2_acc_1725_nl;
  wire[10:0] Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1714_nl;
  wire[11:0] nl_Accum2_acc_1714_nl;
  wire[10:0] Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1727_nl;
  wire[14:0] nl_Accum2_acc_1727_nl;
  wire[11:0] Accum2_acc_1723_nl;
  wire[13:0] nl_Accum2_acc_1723_nl;
  wire[10:0] Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1743_nl;
  wire[14:0] nl_Accum2_acc_1743_nl;
  wire[11:0] Accum2_acc_1740_nl;
  wire[13:0] nl_Accum2_acc_1740_nl;
  wire[10:0] Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1729_nl;
  wire[11:0] nl_Accum2_acc_1729_nl;
  wire[10:0] Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1742_nl;
  wire[14:0] nl_Accum2_acc_1742_nl;
  wire[11:0] Accum2_acc_1738_nl;
  wire[13:0] nl_Accum2_acc_1738_nl;
  wire[10:0] Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1758_nl;
  wire[14:0] nl_Accum2_acc_1758_nl;
  wire[11:0] Accum2_acc_1755_nl;
  wire[13:0] nl_Accum2_acc_1755_nl;
  wire[10:0] Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1744_nl;
  wire[11:0] nl_Accum2_acc_1744_nl;
  wire[10:0] Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1757_nl;
  wire[14:0] nl_Accum2_acc_1757_nl;
  wire[11:0] Accum2_acc_1753_nl;
  wire[13:0] nl_Accum2_acc_1753_nl;
  wire[10:0] Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1773_nl;
  wire[14:0] nl_Accum2_acc_1773_nl;
  wire[11:0] Accum2_acc_1770_nl;
  wire[13:0] nl_Accum2_acc_1770_nl;
  wire[10:0] Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1759_nl;
  wire[11:0] nl_Accum2_acc_1759_nl;
  wire[10:0] Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1772_nl;
  wire[14:0] nl_Accum2_acc_1772_nl;
  wire[11:0] Accum2_acc_1768_nl;
  wire[13:0] nl_Accum2_acc_1768_nl;
  wire[10:0] Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1788_nl;
  wire[14:0] nl_Accum2_acc_1788_nl;
  wire[11:0] Accum2_acc_1785_nl;
  wire[13:0] nl_Accum2_acc_1785_nl;
  wire[10:0] Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1774_nl;
  wire[11:0] nl_Accum2_acc_1774_nl;
  wire[10:0] Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1787_nl;
  wire[14:0] nl_Accum2_acc_1787_nl;
  wire[11:0] Accum2_acc_1783_nl;
  wire[13:0] nl_Accum2_acc_1783_nl;
  wire[10:0] Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1803_nl;
  wire[14:0] nl_Accum2_acc_1803_nl;
  wire[11:0] Accum2_acc_1800_nl;
  wire[13:0] nl_Accum2_acc_1800_nl;
  wire[10:0] Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1789_nl;
  wire[11:0] nl_Accum2_acc_1789_nl;
  wire[10:0] Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1802_nl;
  wire[14:0] nl_Accum2_acc_1802_nl;
  wire[11:0] Accum2_acc_1798_nl;
  wire[13:0] nl_Accum2_acc_1798_nl;
  wire[10:0] Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1818_nl;
  wire[14:0] nl_Accum2_acc_1818_nl;
  wire[11:0] Accum2_acc_1815_nl;
  wire[13:0] nl_Accum2_acc_1815_nl;
  wire[10:0] Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1804_nl;
  wire[11:0] nl_Accum2_acc_1804_nl;
  wire[10:0] Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1817_nl;
  wire[14:0] nl_Accum2_acc_1817_nl;
  wire[11:0] Accum2_acc_1813_nl;
  wire[13:0] nl_Accum2_acc_1813_nl;
  wire[10:0] Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1833_nl;
  wire[14:0] nl_Accum2_acc_1833_nl;
  wire[11:0] Accum2_acc_1830_nl;
  wire[13:0] nl_Accum2_acc_1830_nl;
  wire[10:0] Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1819_nl;
  wire[11:0] nl_Accum2_acc_1819_nl;
  wire[10:0] Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1832_nl;
  wire[14:0] nl_Accum2_acc_1832_nl;
  wire[11:0] Accum2_acc_1828_nl;
  wire[13:0] nl_Accum2_acc_1828_nl;
  wire[10:0] Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1848_nl;
  wire[14:0] nl_Accum2_acc_1848_nl;
  wire[11:0] Accum2_acc_1845_nl;
  wire[13:0] nl_Accum2_acc_1845_nl;
  wire[10:0] Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1834_nl;
  wire[11:0] nl_Accum2_acc_1834_nl;
  wire[10:0] Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1847_nl;
  wire[14:0] nl_Accum2_acc_1847_nl;
  wire[11:0] Accum2_acc_1843_nl;
  wire[13:0] nl_Accum2_acc_1843_nl;
  wire[10:0] Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1863_nl;
  wire[14:0] nl_Accum2_acc_1863_nl;
  wire[11:0] Accum2_acc_1860_nl;
  wire[13:0] nl_Accum2_acc_1860_nl;
  wire[10:0] Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1849_nl;
  wire[11:0] nl_Accum2_acc_1849_nl;
  wire[10:0] Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1862_nl;
  wire[14:0] nl_Accum2_acc_1862_nl;
  wire[11:0] Accum2_acc_1858_nl;
  wire[13:0] nl_Accum2_acc_1858_nl;
  wire[10:0] Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1878_nl;
  wire[14:0] nl_Accum2_acc_1878_nl;
  wire[11:0] Accum2_acc_1875_nl;
  wire[13:0] nl_Accum2_acc_1875_nl;
  wire[10:0] Product1_3_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1864_nl;
  wire[11:0] nl_Accum2_acc_1864_nl;
  wire[10:0] Product1_15_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1877_nl;
  wire[14:0] nl_Accum2_acc_1877_nl;
  wire[11:0] Accum2_acc_1873_nl;
  wire[13:0] nl_Accum2_acc_1873_nl;
  wire[10:0] Product1_11_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1893_nl;
  wire[14:0] nl_Accum2_acc_1893_nl;
  wire[11:0] Accum2_acc_1890_nl;
  wire[13:0] nl_Accum2_acc_1890_nl;
  wire[10:0] Product1_3_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1879_nl;
  wire[11:0] nl_Accum2_acc_1879_nl;
  wire[10:0] Product1_15_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1892_nl;
  wire[14:0] nl_Accum2_acc_1892_nl;
  wire[11:0] Accum2_acc_1888_nl;
  wire[13:0] nl_Accum2_acc_1888_nl;
  wire[10:0] Product1_11_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1908_nl;
  wire[14:0] nl_Accum2_acc_1908_nl;
  wire[11:0] Accum2_acc_1905_nl;
  wire[13:0] nl_Accum2_acc_1905_nl;
  wire[10:0] Product1_3_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1894_nl;
  wire[11:0] nl_Accum2_acc_1894_nl;
  wire[10:0] Product1_15_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1907_nl;
  wire[14:0] nl_Accum2_acc_1907_nl;
  wire[11:0] Accum2_acc_1903_nl;
  wire[13:0] nl_Accum2_acc_1903_nl;
  wire[10:0] Product1_11_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1923_nl;
  wire[14:0] nl_Accum2_acc_1923_nl;
  wire[11:0] Accum2_acc_1920_nl;
  wire[13:0] nl_Accum2_acc_1920_nl;
  wire[10:0] Product1_3_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1909_nl;
  wire[11:0] nl_Accum2_acc_1909_nl;
  wire[10:0] Product1_15_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1922_nl;
  wire[14:0] nl_Accum2_acc_1922_nl;
  wire[11:0] Accum2_acc_1918_nl;
  wire[13:0] nl_Accum2_acc_1918_nl;
  wire[10:0] Product1_11_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1938_nl;
  wire[14:0] nl_Accum2_acc_1938_nl;
  wire[11:0] Accum2_acc_1935_nl;
  wire[13:0] nl_Accum2_acc_1935_nl;
  wire[10:0] Product1_3_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1924_nl;
  wire[11:0] nl_Accum2_acc_1924_nl;
  wire[10:0] Product1_15_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1937_nl;
  wire[14:0] nl_Accum2_acc_1937_nl;
  wire[11:0] Accum2_acc_1933_nl;
  wire[13:0] nl_Accum2_acc_1933_nl;
  wire[10:0] Product1_11_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1953_nl;
  wire[14:0] nl_Accum2_acc_1953_nl;
  wire[11:0] Accum2_acc_1950_nl;
  wire[13:0] nl_Accum2_acc_1950_nl;
  wire[10:0] Product1_3_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_3_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_4_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_4_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_5_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_5_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_6_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_6_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Accum2_acc_1939_nl;
  wire[11:0] nl_Accum2_acc_1939_nl;
  wire[10:0] Product1_15_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_15_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_16_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_16_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_1_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_1_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_2_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_2_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[11:0] Accum2_acc_1952_nl;
  wire[14:0] nl_Accum2_acc_1952_nl;
  wire[11:0] Accum2_acc_1948_nl;
  wire[13:0] nl_Accum2_acc_1948_nl;
  wire[10:0] Product1_11_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_11_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_12_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_12_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_13_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_13_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_14_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_14_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_7_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_7_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_8_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_8_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_9_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_9_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[10:0] Product1_10_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire signed [11:0] nl_Product1_10_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_192_nl;
  wire[6:0] nl_Accum2_1_acc_192_nl;
  wire[14:0] Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_193_nl;
  wire[6:0] nl_Accum2_1_acc_193_nl;
  wire[14:0] Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[5:0] Accum2_1_acc_191_nl;
  wire[6:0] nl_Accum2_1_acc_191_nl;
  wire[14:0] Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[14:0] Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire signed [15:0] nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl;
  wire[12:0] operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl;
  wire[13:0] nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;
  wire[2:0] nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl;

  // Interconnect Declarations for Component Instantiations 
  converterBlock_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd96)) input_1_rsci (
      .dat(input_1_rsc_dat),
      .idat(input_1_rsci_idat)
    );
  converterBlock_ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd2)) layer7_out_rsci (
      .idat(layer7_out_rsci_idat),
      .dat(layer7_out_rsc_dat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd5120)) w2_rsci (
      .dat(w2_rsc_dat),
      .idat(w2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd320)) b2_rsci (
      .dat(b2_rsc_dat),
      .idat(b2_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd960)) w5_rsci (
      .dat(w5_rsc_dat),
      .idat(w5_rsci_idat)
    );
  converterBlock_ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd15)) b5_rsci (
      .dat(b5_rsc_dat),
      .idat(b5_rsci_idat)
    );
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1 = (layer3_out_0_15_4_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[964:960]));
  assign Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1284:1280]));
  assign Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1604:1600]));
  assign Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1924:1920]));
  assign Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1965_nl = conv_s2s_11_12(Product1_4_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_7_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1965_nl = nl_Accum2_acc_1965_nl[11:0];
  assign nl_Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4804:4800]));
  assign Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1954_nl = Product1_16_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[4:0]);
  assign Accum2_acc_1954_nl = nl_Accum2_acc_1954_nl[10:0];
  assign nl_Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[4:0]));
  assign Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[324:320]));
  assign Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[644:640]));
  assign Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1968_nl = Accum2_acc_1965_nl + conv_s2s_11_12(Accum2_acc_1954_nl)
      + conv_s2s_11_12(Product1_1_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_3_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1968_nl = nl_Accum2_acc_1968_nl[11:0];
  assign nl_Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3524:3520]));
  assign Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3844:3840]));
  assign Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4164:4160]));
  assign Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4484:4480]));
  assign Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1963_nl = conv_s2s_11_12(Product1_12_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_15_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1963_nl = nl_Accum2_acc_1963_nl[11:0];
  assign nl_Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2244:2240]));
  assign Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2564:2560]));
  assign Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2884:2880]));
  assign Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3204:3200]));
  assign Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1967_nl = Accum2_acc_1963_nl + conv_s2s_11_12(Product1_8_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_11_Product2_1_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1967_nl = nl_Accum2_acc_1967_nl[11:0];
  assign nl_layer3_out_0_15_4_sva_1 = Accum2_acc_1968_nl + Accum2_acc_1967_nl;
  assign layer3_out_0_15_4_sva_1 = nl_layer3_out_0_15_4_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 = (Accum2_acc_65_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[649:645]));
  assign Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[969:965]));
  assign Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1289:1285]));
  assign Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1609:1605]));
  assign Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1020_nl = conv_s2s_11_12(Product1_3_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1020_nl = nl_Accum2_acc_1020_nl[11:0];
  assign nl_Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4489:4485]));
  assign Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1017_nl = Product1_15_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[9:5]);
  assign Accum2_acc_1017_nl = nl_Accum2_acc_1017_nl[10:0];
  assign nl_Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4809:4805]));
  assign Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[9:5]));
  assign Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[329:325]));
  assign Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_nl = Accum2_acc_1020_nl + conv_s2s_11_12(Accum2_acc_1017_nl)
      + conv_s2s_11_12(Product1_16_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_nl = nl_Accum2_acc_nl[11:0];
  assign nl_Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3209:3205]));
  assign Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3529:3525]));
  assign Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3849:3845]));
  assign Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4169:4165]));
  assign Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1018_nl = conv_s2s_11_12(Product1_11_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1018_nl = nl_Accum2_acc_1018_nl[11:0];
  assign nl_Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1929:1925]));
  assign Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2249:2245]));
  assign Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2569:2565]));
  assign Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2889:2885]));
  assign Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1022_nl = Accum2_acc_1018_nl + conv_s2s_11_12(Product1_7_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_2_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1022_nl = nl_Accum2_acc_1022_nl[11:0];
  assign nl_Accum2_acc_65_psp_sva_1 = Accum2_acc_nl + Accum2_acc_1022_nl;
  assign Accum2_acc_65_psp_sva_1 = nl_Accum2_acc_65_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 = (Accum2_acc_66_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[654:650]));
  assign Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[974:970]));
  assign Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1294:1290]));
  assign Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1614:1610]));
  assign Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1035_nl = conv_s2s_11_12(Product1_3_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1035_nl = nl_Accum2_acc_1035_nl[11:0];
  assign nl_Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4494:4490]));
  assign Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1024_nl = Product1_15_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[14:10]);
  assign Accum2_acc_1024_nl = nl_Accum2_acc_1024_nl[10:0];
  assign nl_Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4814:4810]));
  assign Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[14:10]));
  assign Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[334:330]));
  assign Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1038_nl = Accum2_acc_1035_nl + conv_s2s_11_12(Accum2_acc_1024_nl)
      + conv_s2s_11_12(Product1_16_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1038_nl = nl_Accum2_acc_1038_nl[11:0];
  assign nl_Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3214:3210]));
  assign Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3534:3530]));
  assign Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3854:3850]));
  assign Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4174:4170]));
  assign Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1033_nl = conv_s2s_11_12(Product1_11_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1033_nl = nl_Accum2_acc_1033_nl[11:0];
  assign nl_Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1934:1930]));
  assign Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2254:2250]));
  assign Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2574:2570]));
  assign Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2894:2890]));
  assign Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1037_nl = Accum2_acc_1033_nl + conv_s2s_11_12(Product1_7_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_3_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1037_nl = nl_Accum2_acc_1037_nl[11:0];
  assign nl_Accum2_acc_66_psp_sva_1 = Accum2_acc_1038_nl + Accum2_acc_1037_nl;
  assign Accum2_acc_66_psp_sva_1 = nl_Accum2_acc_66_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 = (Accum2_acc_67_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[659:655]));
  assign Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[979:975]));
  assign Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1299:1295]));
  assign Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1619:1615]));
  assign Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1050_nl = conv_s2s_11_12(Product1_3_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1050_nl = nl_Accum2_acc_1050_nl[11:0];
  assign nl_Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4499:4495]));
  assign Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1039_nl = Product1_15_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[19:15]);
  assign Accum2_acc_1039_nl = nl_Accum2_acc_1039_nl[10:0];
  assign nl_Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4819:4815]));
  assign Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[19:15]));
  assign Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[339:335]));
  assign Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1053_nl = Accum2_acc_1050_nl + conv_s2s_11_12(Accum2_acc_1039_nl)
      + conv_s2s_11_12(Product1_16_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1053_nl = nl_Accum2_acc_1053_nl[11:0];
  assign nl_Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3219:3215]));
  assign Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3539:3535]));
  assign Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3859:3855]));
  assign Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4179:4175]));
  assign Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1048_nl = conv_s2s_11_12(Product1_11_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1048_nl = nl_Accum2_acc_1048_nl[11:0];
  assign nl_Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1939:1935]));
  assign Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2259:2255]));
  assign Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2579:2575]));
  assign Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2899:2895]));
  assign Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1052_nl = Accum2_acc_1048_nl + conv_s2s_11_12(Product1_7_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_4_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1052_nl = nl_Accum2_acc_1052_nl[11:0];
  assign nl_Accum2_acc_67_psp_sva_1 = Accum2_acc_1053_nl + Accum2_acc_1052_nl;
  assign Accum2_acc_67_psp_sva_1 = nl_Accum2_acc_67_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 = (Accum2_acc_68_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[664:660]));
  assign Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[984:980]));
  assign Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1304:1300]));
  assign Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1624:1620]));
  assign Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1065_nl = conv_s2s_11_12(Product1_3_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1065_nl = nl_Accum2_acc_1065_nl[11:0];
  assign nl_Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4504:4500]));
  assign Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1054_nl = Product1_15_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[24:20]);
  assign Accum2_acc_1054_nl = nl_Accum2_acc_1054_nl[10:0];
  assign nl_Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4824:4820]));
  assign Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[24:20]));
  assign Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[344:340]));
  assign Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1068_nl = Accum2_acc_1065_nl + conv_s2s_11_12(Accum2_acc_1054_nl)
      + conv_s2s_11_12(Product1_16_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1068_nl = nl_Accum2_acc_1068_nl[11:0];
  assign nl_Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3224:3220]));
  assign Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3544:3540]));
  assign Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3864:3860]));
  assign Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4184:4180]));
  assign Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1063_nl = conv_s2s_11_12(Product1_11_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1063_nl = nl_Accum2_acc_1063_nl[11:0];
  assign nl_Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1944:1940]));
  assign Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2264:2260]));
  assign Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2584:2580]));
  assign Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2904:2900]));
  assign Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1067_nl = Accum2_acc_1063_nl + conv_s2s_11_12(Product1_7_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_5_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1067_nl = nl_Accum2_acc_1067_nl[11:0];
  assign nl_Accum2_acc_68_psp_sva_1 = Accum2_acc_1068_nl + Accum2_acc_1067_nl;
  assign Accum2_acc_68_psp_sva_1 = nl_Accum2_acc_68_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 = (Accum2_acc_69_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[669:665]));
  assign Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[989:985]));
  assign Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1309:1305]));
  assign Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1629:1625]));
  assign Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1080_nl = conv_s2s_11_12(Product1_3_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1080_nl = nl_Accum2_acc_1080_nl[11:0];
  assign nl_Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4509:4505]));
  assign Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1069_nl = Product1_15_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[29:25]);
  assign Accum2_acc_1069_nl = nl_Accum2_acc_1069_nl[10:0];
  assign nl_Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4829:4825]));
  assign Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[29:25]));
  assign Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[349:345]));
  assign Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1083_nl = Accum2_acc_1080_nl + conv_s2s_11_12(Accum2_acc_1069_nl)
      + conv_s2s_11_12(Product1_16_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1083_nl = nl_Accum2_acc_1083_nl[11:0];
  assign nl_Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3229:3225]));
  assign Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3549:3545]));
  assign Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3869:3865]));
  assign Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4189:4185]));
  assign Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1078_nl = conv_s2s_11_12(Product1_11_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1078_nl = nl_Accum2_acc_1078_nl[11:0];
  assign nl_Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1949:1945]));
  assign Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2269:2265]));
  assign Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2589:2585]));
  assign Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2909:2905]));
  assign Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1082_nl = Accum2_acc_1078_nl + conv_s2s_11_12(Product1_7_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_6_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1082_nl = nl_Accum2_acc_1082_nl[11:0];
  assign nl_Accum2_acc_69_psp_sva_1 = Accum2_acc_1083_nl + Accum2_acc_1082_nl;
  assign Accum2_acc_69_psp_sva_1 = nl_Accum2_acc_69_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 = (Accum2_acc_70_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[674:670]));
  assign Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[994:990]));
  assign Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1314:1310]));
  assign Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1634:1630]));
  assign Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1095_nl = conv_s2s_11_12(Product1_3_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1095_nl = nl_Accum2_acc_1095_nl[11:0];
  assign nl_Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4514:4510]));
  assign Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1084_nl = Product1_15_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[34:30]);
  assign Accum2_acc_1084_nl = nl_Accum2_acc_1084_nl[10:0];
  assign nl_Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4834:4830]));
  assign Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[34:30]));
  assign Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[354:350]));
  assign Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1098_nl = Accum2_acc_1095_nl + conv_s2s_11_12(Accum2_acc_1084_nl)
      + conv_s2s_11_12(Product1_16_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1098_nl = nl_Accum2_acc_1098_nl[11:0];
  assign nl_Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3234:3230]));
  assign Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3554:3550]));
  assign Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3874:3870]));
  assign Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4194:4190]));
  assign Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1093_nl = conv_s2s_11_12(Product1_11_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1093_nl = nl_Accum2_acc_1093_nl[11:0];
  assign nl_Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1954:1950]));
  assign Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2274:2270]));
  assign Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2594:2590]));
  assign Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2914:2910]));
  assign Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1097_nl = Accum2_acc_1093_nl + conv_s2s_11_12(Product1_7_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_7_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1097_nl = nl_Accum2_acc_1097_nl[11:0];
  assign nl_Accum2_acc_70_psp_sva_1 = Accum2_acc_1098_nl + Accum2_acc_1097_nl;
  assign Accum2_acc_70_psp_sva_1 = nl_Accum2_acc_70_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 = (Accum2_acc_71_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[679:675]));
  assign Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[999:995]));
  assign Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1319:1315]));
  assign Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1639:1635]));
  assign Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1110_nl = conv_s2s_11_12(Product1_3_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1110_nl = nl_Accum2_acc_1110_nl[11:0];
  assign nl_Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4519:4515]));
  assign Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1099_nl = Product1_15_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[39:35]);
  assign Accum2_acc_1099_nl = nl_Accum2_acc_1099_nl[10:0];
  assign nl_Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4839:4835]));
  assign Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[39:35]));
  assign Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[359:355]));
  assign Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1113_nl = Accum2_acc_1110_nl + conv_s2s_11_12(Accum2_acc_1099_nl)
      + conv_s2s_11_12(Product1_16_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1113_nl = nl_Accum2_acc_1113_nl[11:0];
  assign nl_Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3239:3235]));
  assign Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3559:3555]));
  assign Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3879:3875]));
  assign Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4199:4195]));
  assign Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1108_nl = conv_s2s_11_12(Product1_11_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1108_nl = nl_Accum2_acc_1108_nl[11:0];
  assign nl_Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1959:1955]));
  assign Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2279:2275]));
  assign Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2599:2595]));
  assign Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2919:2915]));
  assign Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1112_nl = Accum2_acc_1108_nl + conv_s2s_11_12(Product1_7_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_8_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1112_nl = nl_Accum2_acc_1112_nl[11:0];
  assign nl_Accum2_acc_71_psp_sva_1 = Accum2_acc_1113_nl + Accum2_acc_1112_nl;
  assign Accum2_acc_71_psp_sva_1 = nl_Accum2_acc_71_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 = (Accum2_acc_72_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[684:680]));
  assign Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1004:1000]));
  assign Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1324:1320]));
  assign Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1644:1640]));
  assign Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1125_nl = conv_s2s_11_12(Product1_3_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1125_nl = nl_Accum2_acc_1125_nl[11:0];
  assign nl_Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4524:4520]));
  assign Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1114_nl = Product1_15_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[44:40]);
  assign Accum2_acc_1114_nl = nl_Accum2_acc_1114_nl[10:0];
  assign nl_Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4844:4840]));
  assign Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[44:40]));
  assign Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[364:360]));
  assign Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1128_nl = Accum2_acc_1125_nl + conv_s2s_11_12(Accum2_acc_1114_nl)
      + conv_s2s_11_12(Product1_16_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1128_nl = nl_Accum2_acc_1128_nl[11:0];
  assign nl_Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3244:3240]));
  assign Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3564:3560]));
  assign Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3884:3880]));
  assign Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4204:4200]));
  assign Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1123_nl = conv_s2s_11_12(Product1_11_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1123_nl = nl_Accum2_acc_1123_nl[11:0];
  assign nl_Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1964:1960]));
  assign Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2284:2280]));
  assign Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2604:2600]));
  assign Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2924:2920]));
  assign Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1127_nl = Accum2_acc_1123_nl + conv_s2s_11_12(Product1_7_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_9_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1127_nl = nl_Accum2_acc_1127_nl[11:0];
  assign nl_Accum2_acc_72_psp_sva_1 = Accum2_acc_1128_nl + Accum2_acc_1127_nl;
  assign Accum2_acc_72_psp_sva_1 = nl_Accum2_acc_72_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 = (Accum2_acc_73_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[689:685]));
  assign Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1009:1005]));
  assign Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1329:1325]));
  assign Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1649:1645]));
  assign Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1140_nl = conv_s2s_11_12(Product1_3_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1140_nl = nl_Accum2_acc_1140_nl[11:0];
  assign nl_Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4529:4525]));
  assign Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1129_nl = Product1_15_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[49:45]);
  assign Accum2_acc_1129_nl = nl_Accum2_acc_1129_nl[10:0];
  assign nl_Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4849:4845]));
  assign Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[49:45]));
  assign Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[369:365]));
  assign Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1143_nl = Accum2_acc_1140_nl + conv_s2s_11_12(Accum2_acc_1129_nl)
      + conv_s2s_11_12(Product1_16_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1143_nl = nl_Accum2_acc_1143_nl[11:0];
  assign nl_Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3249:3245]));
  assign Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3569:3565]));
  assign Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3889:3885]));
  assign Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4209:4205]));
  assign Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1138_nl = conv_s2s_11_12(Product1_11_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1138_nl = nl_Accum2_acc_1138_nl[11:0];
  assign nl_Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1969:1965]));
  assign Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2289:2285]));
  assign Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2609:2605]));
  assign Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2929:2925]));
  assign Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1142_nl = Accum2_acc_1138_nl + conv_s2s_11_12(Product1_7_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_10_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1142_nl = nl_Accum2_acc_1142_nl[11:0];
  assign nl_Accum2_acc_73_psp_sva_1 = Accum2_acc_1143_nl + Accum2_acc_1142_nl;
  assign Accum2_acc_73_psp_sva_1 = nl_Accum2_acc_73_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 = (Accum2_acc_74_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[694:690]));
  assign Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1014:1010]));
  assign Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1334:1330]));
  assign Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1654:1650]));
  assign Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1155_nl = conv_s2s_11_12(Product1_3_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1155_nl = nl_Accum2_acc_1155_nl[11:0];
  assign nl_Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4534:4530]));
  assign Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1144_nl = Product1_15_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[54:50]);
  assign Accum2_acc_1144_nl = nl_Accum2_acc_1144_nl[10:0];
  assign nl_Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4854:4850]));
  assign Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[54:50]));
  assign Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[374:370]));
  assign Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1158_nl = Accum2_acc_1155_nl + conv_s2s_11_12(Accum2_acc_1144_nl)
      + conv_s2s_11_12(Product1_16_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1158_nl = nl_Accum2_acc_1158_nl[11:0];
  assign nl_Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3254:3250]));
  assign Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3574:3570]));
  assign Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3894:3890]));
  assign Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4214:4210]));
  assign Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1153_nl = conv_s2s_11_12(Product1_11_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1153_nl = nl_Accum2_acc_1153_nl[11:0];
  assign nl_Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1974:1970]));
  assign Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2294:2290]));
  assign Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2614:2610]));
  assign Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2934:2930]));
  assign Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1157_nl = Accum2_acc_1153_nl + conv_s2s_11_12(Product1_7_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_11_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1157_nl = nl_Accum2_acc_1157_nl[11:0];
  assign nl_Accum2_acc_74_psp_sva_1 = Accum2_acc_1158_nl + Accum2_acc_1157_nl;
  assign Accum2_acc_74_psp_sva_1 = nl_Accum2_acc_74_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 = (Accum2_acc_75_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[699:695]));
  assign Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1019:1015]));
  assign Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1339:1335]));
  assign Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1659:1655]));
  assign Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1170_nl = conv_s2s_11_12(Product1_3_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1170_nl = nl_Accum2_acc_1170_nl[11:0];
  assign nl_Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4539:4535]));
  assign Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1159_nl = Product1_15_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[59:55]);
  assign Accum2_acc_1159_nl = nl_Accum2_acc_1159_nl[10:0];
  assign nl_Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4859:4855]));
  assign Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[59:55]));
  assign Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[379:375]));
  assign Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1173_nl = Accum2_acc_1170_nl + conv_s2s_11_12(Accum2_acc_1159_nl)
      + conv_s2s_11_12(Product1_16_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1173_nl = nl_Accum2_acc_1173_nl[11:0];
  assign nl_Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3259:3255]));
  assign Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3579:3575]));
  assign Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3899:3895]));
  assign Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4219:4215]));
  assign Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1168_nl = conv_s2s_11_12(Product1_11_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1168_nl = nl_Accum2_acc_1168_nl[11:0];
  assign nl_Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1979:1975]));
  assign Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2299:2295]));
  assign Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2619:2615]));
  assign Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2939:2935]));
  assign Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1172_nl = Accum2_acc_1168_nl + conv_s2s_11_12(Product1_7_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_12_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1172_nl = nl_Accum2_acc_1172_nl[11:0];
  assign nl_Accum2_acc_75_psp_sva_1 = Accum2_acc_1173_nl + Accum2_acc_1172_nl;
  assign Accum2_acc_75_psp_sva_1 = nl_Accum2_acc_75_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 = (Accum2_acc_76_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[704:700]));
  assign Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1024:1020]));
  assign Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1344:1340]));
  assign Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1664:1660]));
  assign Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1185_nl = conv_s2s_11_12(Product1_3_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1185_nl = nl_Accum2_acc_1185_nl[11:0];
  assign nl_Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4544:4540]));
  assign Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1174_nl = Product1_15_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[64:60]);
  assign Accum2_acc_1174_nl = nl_Accum2_acc_1174_nl[10:0];
  assign nl_Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4864:4860]));
  assign Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[64:60]));
  assign Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[384:380]));
  assign Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1188_nl = Accum2_acc_1185_nl + conv_s2s_11_12(Accum2_acc_1174_nl)
      + conv_s2s_11_12(Product1_16_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1188_nl = nl_Accum2_acc_1188_nl[11:0];
  assign nl_Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3264:3260]));
  assign Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3584:3580]));
  assign Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3904:3900]));
  assign Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4224:4220]));
  assign Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1183_nl = conv_s2s_11_12(Product1_11_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1183_nl = nl_Accum2_acc_1183_nl[11:0];
  assign nl_Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1984:1980]));
  assign Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2304:2300]));
  assign Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2624:2620]));
  assign Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2944:2940]));
  assign Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1187_nl = Accum2_acc_1183_nl + conv_s2s_11_12(Product1_7_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_13_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1187_nl = nl_Accum2_acc_1187_nl[11:0];
  assign nl_Accum2_acc_76_psp_sva_1 = Accum2_acc_1188_nl + Accum2_acc_1187_nl;
  assign Accum2_acc_76_psp_sva_1 = nl_Accum2_acc_76_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 = (Accum2_acc_77_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[709:705]));
  assign Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1029:1025]));
  assign Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1349:1345]));
  assign Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1669:1665]));
  assign Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1200_nl = conv_s2s_11_12(Product1_3_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1200_nl = nl_Accum2_acc_1200_nl[11:0];
  assign nl_Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4549:4545]));
  assign Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1189_nl = Product1_15_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[69:65]);
  assign Accum2_acc_1189_nl = nl_Accum2_acc_1189_nl[10:0];
  assign nl_Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4869:4865]));
  assign Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[69:65]));
  assign Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[389:385]));
  assign Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1203_nl = Accum2_acc_1200_nl + conv_s2s_11_12(Accum2_acc_1189_nl)
      + conv_s2s_11_12(Product1_16_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1203_nl = nl_Accum2_acc_1203_nl[11:0];
  assign nl_Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3269:3265]));
  assign Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3589:3585]));
  assign Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3909:3905]));
  assign Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4229:4225]));
  assign Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1198_nl = conv_s2s_11_12(Product1_11_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1198_nl = nl_Accum2_acc_1198_nl[11:0];
  assign nl_Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1989:1985]));
  assign Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2309:2305]));
  assign Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2629:2625]));
  assign Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2949:2945]));
  assign Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1202_nl = Accum2_acc_1198_nl + conv_s2s_11_12(Product1_7_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_14_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1202_nl = nl_Accum2_acc_1202_nl[11:0];
  assign nl_Accum2_acc_77_psp_sva_1 = Accum2_acc_1203_nl + Accum2_acc_1202_nl;
  assign Accum2_acc_77_psp_sva_1 = nl_Accum2_acc_77_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 = (Accum2_acc_78_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[714:710]));
  assign Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1034:1030]));
  assign Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1354:1350]));
  assign Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1674:1670]));
  assign Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1215_nl = conv_s2s_11_12(Product1_3_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1215_nl = nl_Accum2_acc_1215_nl[11:0];
  assign nl_Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4554:4550]));
  assign Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1204_nl = Product1_15_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[74:70]);
  assign Accum2_acc_1204_nl = nl_Accum2_acc_1204_nl[10:0];
  assign nl_Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4874:4870]));
  assign Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[74:70]));
  assign Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[394:390]));
  assign Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1218_nl = Accum2_acc_1215_nl + conv_s2s_11_12(Accum2_acc_1204_nl)
      + conv_s2s_11_12(Product1_16_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1218_nl = nl_Accum2_acc_1218_nl[11:0];
  assign nl_Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3274:3270]));
  assign Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3594:3590]));
  assign Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3914:3910]));
  assign Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4234:4230]));
  assign Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1213_nl = conv_s2s_11_12(Product1_11_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1213_nl = nl_Accum2_acc_1213_nl[11:0];
  assign nl_Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1994:1990]));
  assign Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2314:2310]));
  assign Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2634:2630]));
  assign Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2954:2950]));
  assign Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1217_nl = Accum2_acc_1213_nl + conv_s2s_11_12(Product1_7_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_15_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1217_nl = nl_Accum2_acc_1217_nl[11:0];
  assign nl_Accum2_acc_78_psp_sva_1 = Accum2_acc_1218_nl + Accum2_acc_1217_nl;
  assign Accum2_acc_78_psp_sva_1 = nl_Accum2_acc_78_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 = (Accum2_acc_79_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[719:715]));
  assign Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1039:1035]));
  assign Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1359:1355]));
  assign Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1679:1675]));
  assign Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1230_nl = conv_s2s_11_12(Product1_3_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1230_nl = nl_Accum2_acc_1230_nl[11:0];
  assign nl_Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4559:4555]));
  assign Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1219_nl = Product1_15_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[79:75]);
  assign Accum2_acc_1219_nl = nl_Accum2_acc_1219_nl[10:0];
  assign nl_Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4879:4875]));
  assign Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[79:75]));
  assign Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[399:395]));
  assign Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1233_nl = Accum2_acc_1230_nl + conv_s2s_11_12(Accum2_acc_1219_nl)
      + conv_s2s_11_12(Product1_16_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1233_nl = nl_Accum2_acc_1233_nl[11:0];
  assign nl_Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3279:3275]));
  assign Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3599:3595]));
  assign Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3919:3915]));
  assign Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4239:4235]));
  assign Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1228_nl = conv_s2s_11_12(Product1_11_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1228_nl = nl_Accum2_acc_1228_nl[11:0];
  assign nl_Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[1999:1995]));
  assign Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2319:2315]));
  assign Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2639:2635]));
  assign Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2959:2955]));
  assign Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1232_nl = Accum2_acc_1228_nl + conv_s2s_11_12(Product1_7_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_16_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1232_nl = nl_Accum2_acc_1232_nl[11:0];
  assign nl_Accum2_acc_79_psp_sva_1 = Accum2_acc_1233_nl + Accum2_acc_1232_nl;
  assign Accum2_acc_79_psp_sva_1 = nl_Accum2_acc_79_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 = (Accum2_acc_80_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[724:720]));
  assign Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1044:1040]));
  assign Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1364:1360]));
  assign Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1684:1680]));
  assign Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1245_nl = conv_s2s_11_12(Product1_3_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1245_nl = nl_Accum2_acc_1245_nl[11:0];
  assign nl_Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4564:4560]));
  assign Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1234_nl = Product1_15_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[84:80]);
  assign Accum2_acc_1234_nl = nl_Accum2_acc_1234_nl[10:0];
  assign nl_Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4884:4880]));
  assign Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[84:80]));
  assign Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[404:400]));
  assign Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1248_nl = Accum2_acc_1245_nl + conv_s2s_11_12(Accum2_acc_1234_nl)
      + conv_s2s_11_12(Product1_16_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1248_nl = nl_Accum2_acc_1248_nl[11:0];
  assign nl_Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3284:3280]));
  assign Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3604:3600]));
  assign Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3924:3920]));
  assign Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4244:4240]));
  assign Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1243_nl = conv_s2s_11_12(Product1_11_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1243_nl = nl_Accum2_acc_1243_nl[11:0];
  assign nl_Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2004:2000]));
  assign Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2324:2320]));
  assign Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2644:2640]));
  assign Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2964:2960]));
  assign Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1247_nl = Accum2_acc_1243_nl + conv_s2s_11_12(Product1_7_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_17_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1247_nl = nl_Accum2_acc_1247_nl[11:0];
  assign nl_Accum2_acc_80_psp_sva_1 = Accum2_acc_1248_nl + Accum2_acc_1247_nl;
  assign Accum2_acc_80_psp_sva_1 = nl_Accum2_acc_80_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 = (Accum2_acc_81_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[729:725]));
  assign Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1049:1045]));
  assign Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1369:1365]));
  assign Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1689:1685]));
  assign Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1260_nl = conv_s2s_11_12(Product1_3_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1260_nl = nl_Accum2_acc_1260_nl[11:0];
  assign nl_Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4569:4565]));
  assign Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1249_nl = Product1_15_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[89:85]);
  assign Accum2_acc_1249_nl = nl_Accum2_acc_1249_nl[10:0];
  assign nl_Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4889:4885]));
  assign Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[89:85]));
  assign Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[409:405]));
  assign Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1263_nl = Accum2_acc_1260_nl + conv_s2s_11_12(Accum2_acc_1249_nl)
      + conv_s2s_11_12(Product1_16_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1263_nl = nl_Accum2_acc_1263_nl[11:0];
  assign nl_Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3289:3285]));
  assign Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3609:3605]));
  assign Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3929:3925]));
  assign Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4249:4245]));
  assign Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1258_nl = conv_s2s_11_12(Product1_11_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1258_nl = nl_Accum2_acc_1258_nl[11:0];
  assign nl_Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2009:2005]));
  assign Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2329:2325]));
  assign Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2649:2645]));
  assign Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2969:2965]));
  assign Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1262_nl = Accum2_acc_1258_nl + conv_s2s_11_12(Product1_7_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_18_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1262_nl = nl_Accum2_acc_1262_nl[11:0];
  assign nl_Accum2_acc_81_psp_sva_1 = Accum2_acc_1263_nl + Accum2_acc_1262_nl;
  assign Accum2_acc_81_psp_sva_1 = nl_Accum2_acc_81_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 = (Accum2_acc_82_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[734:730]));
  assign Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1054:1050]));
  assign Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1374:1370]));
  assign Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1694:1690]));
  assign Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1275_nl = conv_s2s_11_12(Product1_3_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1275_nl = nl_Accum2_acc_1275_nl[11:0];
  assign nl_Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4574:4570]));
  assign Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1264_nl = Product1_15_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[94:90]);
  assign Accum2_acc_1264_nl = nl_Accum2_acc_1264_nl[10:0];
  assign nl_Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4894:4890]));
  assign Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[94:90]));
  assign Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[414:410]));
  assign Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1278_nl = Accum2_acc_1275_nl + conv_s2s_11_12(Accum2_acc_1264_nl)
      + conv_s2s_11_12(Product1_16_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1278_nl = nl_Accum2_acc_1278_nl[11:0];
  assign nl_Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3294:3290]));
  assign Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3614:3610]));
  assign Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3934:3930]));
  assign Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4254:4250]));
  assign Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1273_nl = conv_s2s_11_12(Product1_11_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1273_nl = nl_Accum2_acc_1273_nl[11:0];
  assign nl_Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2014:2010]));
  assign Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2334:2330]));
  assign Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2654:2650]));
  assign Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2974:2970]));
  assign Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1277_nl = Accum2_acc_1273_nl + conv_s2s_11_12(Product1_7_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_19_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1277_nl = nl_Accum2_acc_1277_nl[11:0];
  assign nl_Accum2_acc_82_psp_sva_1 = Accum2_acc_1278_nl + Accum2_acc_1277_nl;
  assign Accum2_acc_82_psp_sva_1 = nl_Accum2_acc_82_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 = (Accum2_acc_83_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[739:735]));
  assign Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1059:1055]));
  assign Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1379:1375]));
  assign Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1699:1695]));
  assign Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1290_nl = conv_s2s_11_12(Product1_3_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1290_nl = nl_Accum2_acc_1290_nl[11:0];
  assign nl_Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4579:4575]));
  assign Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1279_nl = Product1_15_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[99:95]);
  assign Accum2_acc_1279_nl = nl_Accum2_acc_1279_nl[10:0];
  assign nl_Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4899:4895]));
  assign Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[99:95]));
  assign Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[419:415]));
  assign Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1293_nl = Accum2_acc_1290_nl + conv_s2s_11_12(Accum2_acc_1279_nl)
      + conv_s2s_11_12(Product1_16_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1293_nl = nl_Accum2_acc_1293_nl[11:0];
  assign nl_Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3299:3295]));
  assign Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3619:3615]));
  assign Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3939:3935]));
  assign Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4259:4255]));
  assign Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1288_nl = conv_s2s_11_12(Product1_11_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1288_nl = nl_Accum2_acc_1288_nl[11:0];
  assign nl_Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2019:2015]));
  assign Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2339:2335]));
  assign Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2659:2655]));
  assign Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2979:2975]));
  assign Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1292_nl = Accum2_acc_1288_nl + conv_s2s_11_12(Product1_7_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_20_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1292_nl = nl_Accum2_acc_1292_nl[11:0];
  assign nl_Accum2_acc_83_psp_sva_1 = Accum2_acc_1293_nl + Accum2_acc_1292_nl;
  assign Accum2_acc_83_psp_sva_1 = nl_Accum2_acc_83_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 = (Accum2_acc_84_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[744:740]));
  assign Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1064:1060]));
  assign Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1384:1380]));
  assign Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1704:1700]));
  assign Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1305_nl = conv_s2s_11_12(Product1_3_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1305_nl = nl_Accum2_acc_1305_nl[11:0];
  assign nl_Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4584:4580]));
  assign Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1294_nl = Product1_15_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[104:100]);
  assign Accum2_acc_1294_nl = nl_Accum2_acc_1294_nl[10:0];
  assign nl_Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4904:4900]));
  assign Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[104:100]));
  assign Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[424:420]));
  assign Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1308_nl = Accum2_acc_1305_nl + conv_s2s_11_12(Accum2_acc_1294_nl)
      + conv_s2s_11_12(Product1_16_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1308_nl = nl_Accum2_acc_1308_nl[11:0];
  assign nl_Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3304:3300]));
  assign Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3624:3620]));
  assign Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3944:3940]));
  assign Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4264:4260]));
  assign Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1303_nl = conv_s2s_11_12(Product1_11_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1303_nl = nl_Accum2_acc_1303_nl[11:0];
  assign nl_Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2024:2020]));
  assign Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2344:2340]));
  assign Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2664:2660]));
  assign Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2984:2980]));
  assign Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1307_nl = Accum2_acc_1303_nl + conv_s2s_11_12(Product1_7_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_21_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1307_nl = nl_Accum2_acc_1307_nl[11:0];
  assign nl_Accum2_acc_84_psp_sva_1 = Accum2_acc_1308_nl + Accum2_acc_1307_nl;
  assign Accum2_acc_84_psp_sva_1 = nl_Accum2_acc_84_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 = (Accum2_acc_85_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[749:745]));
  assign Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1069:1065]));
  assign Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1389:1385]));
  assign Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1709:1705]));
  assign Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1320_nl = conv_s2s_11_12(Product1_3_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1320_nl = nl_Accum2_acc_1320_nl[11:0];
  assign nl_Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4589:4585]));
  assign Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1309_nl = Product1_15_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[109:105]);
  assign Accum2_acc_1309_nl = nl_Accum2_acc_1309_nl[10:0];
  assign nl_Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4909:4905]));
  assign Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[109:105]));
  assign Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[429:425]));
  assign Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1323_nl = Accum2_acc_1320_nl + conv_s2s_11_12(Accum2_acc_1309_nl)
      + conv_s2s_11_12(Product1_16_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1323_nl = nl_Accum2_acc_1323_nl[11:0];
  assign nl_Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3309:3305]));
  assign Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3629:3625]));
  assign Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3949:3945]));
  assign Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4269:4265]));
  assign Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1318_nl = conv_s2s_11_12(Product1_11_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1318_nl = nl_Accum2_acc_1318_nl[11:0];
  assign nl_Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2029:2025]));
  assign Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2349:2345]));
  assign Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2669:2665]));
  assign Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2989:2985]));
  assign Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1322_nl = Accum2_acc_1318_nl + conv_s2s_11_12(Product1_7_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_22_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1322_nl = nl_Accum2_acc_1322_nl[11:0];
  assign nl_Accum2_acc_85_psp_sva_1 = Accum2_acc_1323_nl + Accum2_acc_1322_nl;
  assign Accum2_acc_85_psp_sva_1 = nl_Accum2_acc_85_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 = (Accum2_acc_86_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[754:750]));
  assign Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1074:1070]));
  assign Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1394:1390]));
  assign Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1714:1710]));
  assign Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1335_nl = conv_s2s_11_12(Product1_3_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1335_nl = nl_Accum2_acc_1335_nl[11:0];
  assign nl_Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4594:4590]));
  assign Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1324_nl = Product1_15_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[114:110]);
  assign Accum2_acc_1324_nl = nl_Accum2_acc_1324_nl[10:0];
  assign nl_Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4914:4910]));
  assign Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[114:110]));
  assign Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[434:430]));
  assign Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1338_nl = Accum2_acc_1335_nl + conv_s2s_11_12(Accum2_acc_1324_nl)
      + conv_s2s_11_12(Product1_16_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1338_nl = nl_Accum2_acc_1338_nl[11:0];
  assign nl_Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3314:3310]));
  assign Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3634:3630]));
  assign Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3954:3950]));
  assign Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4274:4270]));
  assign Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1333_nl = conv_s2s_11_12(Product1_11_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1333_nl = nl_Accum2_acc_1333_nl[11:0];
  assign nl_Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2034:2030]));
  assign Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2354:2350]));
  assign Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2674:2670]));
  assign Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2994:2990]));
  assign Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1337_nl = Accum2_acc_1333_nl + conv_s2s_11_12(Product1_7_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_23_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1337_nl = nl_Accum2_acc_1337_nl[11:0];
  assign nl_Accum2_acc_86_psp_sva_1 = Accum2_acc_1338_nl + Accum2_acc_1337_nl;
  assign Accum2_acc_86_psp_sva_1 = nl_Accum2_acc_86_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 = (Accum2_acc_87_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[759:755]));
  assign Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1079:1075]));
  assign Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1399:1395]));
  assign Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1719:1715]));
  assign Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1350_nl = conv_s2s_11_12(Product1_3_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1350_nl = nl_Accum2_acc_1350_nl[11:0];
  assign nl_Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4599:4595]));
  assign Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1339_nl = Product1_15_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[119:115]);
  assign Accum2_acc_1339_nl = nl_Accum2_acc_1339_nl[10:0];
  assign nl_Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4919:4915]));
  assign Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[119:115]));
  assign Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[439:435]));
  assign Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1353_nl = Accum2_acc_1350_nl + conv_s2s_11_12(Accum2_acc_1339_nl)
      + conv_s2s_11_12(Product1_16_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1353_nl = nl_Accum2_acc_1353_nl[11:0];
  assign nl_Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3319:3315]));
  assign Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3639:3635]));
  assign Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3959:3955]));
  assign Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4279:4275]));
  assign Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1348_nl = conv_s2s_11_12(Product1_11_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1348_nl = nl_Accum2_acc_1348_nl[11:0];
  assign nl_Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2039:2035]));
  assign Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2359:2355]));
  assign Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2679:2675]));
  assign Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[2999:2995]));
  assign Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1352_nl = Accum2_acc_1348_nl + conv_s2s_11_12(Product1_7_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_24_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1352_nl = nl_Accum2_acc_1352_nl[11:0];
  assign nl_Accum2_acc_87_psp_sva_1 = Accum2_acc_1353_nl + Accum2_acc_1352_nl;
  assign Accum2_acc_87_psp_sva_1 = nl_Accum2_acc_87_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 = (Accum2_acc_88_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[764:760]));
  assign Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1084:1080]));
  assign Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1404:1400]));
  assign Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1724:1720]));
  assign Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1365_nl = conv_s2s_11_12(Product1_3_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1365_nl = nl_Accum2_acc_1365_nl[11:0];
  assign nl_Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4604:4600]));
  assign Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1354_nl = Product1_15_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[124:120]);
  assign Accum2_acc_1354_nl = nl_Accum2_acc_1354_nl[10:0];
  assign nl_Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4924:4920]));
  assign Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[124:120]));
  assign Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[444:440]));
  assign Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1368_nl = Accum2_acc_1365_nl + conv_s2s_11_12(Accum2_acc_1354_nl)
      + conv_s2s_11_12(Product1_16_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1368_nl = nl_Accum2_acc_1368_nl[11:0];
  assign nl_Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3324:3320]));
  assign Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3644:3640]));
  assign Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3964:3960]));
  assign Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4284:4280]));
  assign Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1363_nl = conv_s2s_11_12(Product1_11_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1363_nl = nl_Accum2_acc_1363_nl[11:0];
  assign nl_Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2044:2040]));
  assign Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2364:2360]));
  assign Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2684:2680]));
  assign Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3004:3000]));
  assign Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1367_nl = Accum2_acc_1363_nl + conv_s2s_11_12(Product1_7_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_25_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1367_nl = nl_Accum2_acc_1367_nl[11:0];
  assign nl_Accum2_acc_88_psp_sva_1 = Accum2_acc_1368_nl + Accum2_acc_1367_nl;
  assign Accum2_acc_88_psp_sva_1 = nl_Accum2_acc_88_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 = (Accum2_acc_89_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[769:765]));
  assign Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1089:1085]));
  assign Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1409:1405]));
  assign Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1729:1725]));
  assign Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1380_nl = conv_s2s_11_12(Product1_3_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1380_nl = nl_Accum2_acc_1380_nl[11:0];
  assign nl_Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4609:4605]));
  assign Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1369_nl = Product1_15_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[129:125]);
  assign Accum2_acc_1369_nl = nl_Accum2_acc_1369_nl[10:0];
  assign nl_Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4929:4925]));
  assign Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[129:125]));
  assign Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[449:445]));
  assign Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1383_nl = Accum2_acc_1380_nl + conv_s2s_11_12(Accum2_acc_1369_nl)
      + conv_s2s_11_12(Product1_16_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1383_nl = nl_Accum2_acc_1383_nl[11:0];
  assign nl_Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3329:3325]));
  assign Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3649:3645]));
  assign Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3969:3965]));
  assign Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4289:4285]));
  assign Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1378_nl = conv_s2s_11_12(Product1_11_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1378_nl = nl_Accum2_acc_1378_nl[11:0];
  assign nl_Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2049:2045]));
  assign Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2369:2365]));
  assign Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2689:2685]));
  assign Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3009:3005]));
  assign Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1382_nl = Accum2_acc_1378_nl + conv_s2s_11_12(Product1_7_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_26_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1382_nl = nl_Accum2_acc_1382_nl[11:0];
  assign nl_Accum2_acc_89_psp_sva_1 = Accum2_acc_1383_nl + Accum2_acc_1382_nl;
  assign Accum2_acc_89_psp_sva_1 = nl_Accum2_acc_89_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 = (Accum2_acc_90_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[774:770]));
  assign Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1094:1090]));
  assign Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1414:1410]));
  assign Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1734:1730]));
  assign Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1395_nl = conv_s2s_11_12(Product1_3_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1395_nl = nl_Accum2_acc_1395_nl[11:0];
  assign nl_Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4614:4610]));
  assign Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1384_nl = Product1_15_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[134:130]);
  assign Accum2_acc_1384_nl = nl_Accum2_acc_1384_nl[10:0];
  assign nl_Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4934:4930]));
  assign Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[134:130]));
  assign Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[454:450]));
  assign Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1398_nl = Accum2_acc_1395_nl + conv_s2s_11_12(Accum2_acc_1384_nl)
      + conv_s2s_11_12(Product1_16_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1398_nl = nl_Accum2_acc_1398_nl[11:0];
  assign nl_Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3334:3330]));
  assign Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3654:3650]));
  assign Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3974:3970]));
  assign Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4294:4290]));
  assign Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1393_nl = conv_s2s_11_12(Product1_11_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1393_nl = nl_Accum2_acc_1393_nl[11:0];
  assign nl_Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2054:2050]));
  assign Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2374:2370]));
  assign Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2694:2690]));
  assign Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3014:3010]));
  assign Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1397_nl = Accum2_acc_1393_nl + conv_s2s_11_12(Product1_7_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_27_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1397_nl = nl_Accum2_acc_1397_nl[11:0];
  assign nl_Accum2_acc_90_psp_sva_1 = Accum2_acc_1398_nl + Accum2_acc_1397_nl;
  assign Accum2_acc_90_psp_sva_1 = nl_Accum2_acc_90_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 = (Accum2_acc_91_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[779:775]));
  assign Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1099:1095]));
  assign Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1419:1415]));
  assign Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1739:1735]));
  assign Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1410_nl = conv_s2s_11_12(Product1_3_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1410_nl = nl_Accum2_acc_1410_nl[11:0];
  assign nl_Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4619:4615]));
  assign Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1399_nl = Product1_15_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[139:135]);
  assign Accum2_acc_1399_nl = nl_Accum2_acc_1399_nl[10:0];
  assign nl_Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4939:4935]));
  assign Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[139:135]));
  assign Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[459:455]));
  assign Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1413_nl = Accum2_acc_1410_nl + conv_s2s_11_12(Accum2_acc_1399_nl)
      + conv_s2s_11_12(Product1_16_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1413_nl = nl_Accum2_acc_1413_nl[11:0];
  assign nl_Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3339:3335]));
  assign Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3659:3655]));
  assign Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3979:3975]));
  assign Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4299:4295]));
  assign Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1408_nl = conv_s2s_11_12(Product1_11_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1408_nl = nl_Accum2_acc_1408_nl[11:0];
  assign nl_Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2059:2055]));
  assign Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2379:2375]));
  assign Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2699:2695]));
  assign Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3019:3015]));
  assign Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1412_nl = Accum2_acc_1408_nl + conv_s2s_11_12(Product1_7_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_28_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1412_nl = nl_Accum2_acc_1412_nl[11:0];
  assign nl_Accum2_acc_91_psp_sva_1 = Accum2_acc_1413_nl + Accum2_acc_1412_nl;
  assign Accum2_acc_91_psp_sva_1 = nl_Accum2_acc_91_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 = (Accum2_acc_92_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[784:780]));
  assign Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1104:1100]));
  assign Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1424:1420]));
  assign Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1744:1740]));
  assign Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1425_nl = conv_s2s_11_12(Product1_3_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1425_nl = nl_Accum2_acc_1425_nl[11:0];
  assign nl_Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4624:4620]));
  assign Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1414_nl = Product1_15_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[144:140]);
  assign Accum2_acc_1414_nl = nl_Accum2_acc_1414_nl[10:0];
  assign nl_Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4944:4940]));
  assign Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[144:140]));
  assign Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[464:460]));
  assign Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1428_nl = Accum2_acc_1425_nl + conv_s2s_11_12(Accum2_acc_1414_nl)
      + conv_s2s_11_12(Product1_16_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1428_nl = nl_Accum2_acc_1428_nl[11:0];
  assign nl_Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3344:3340]));
  assign Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3664:3660]));
  assign Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3984:3980]));
  assign Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4304:4300]));
  assign Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1423_nl = conv_s2s_11_12(Product1_11_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1423_nl = nl_Accum2_acc_1423_nl[11:0];
  assign nl_Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2064:2060]));
  assign Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2384:2380]));
  assign Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2704:2700]));
  assign Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3024:3020]));
  assign Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1427_nl = Accum2_acc_1423_nl + conv_s2s_11_12(Product1_7_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_29_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1427_nl = nl_Accum2_acc_1427_nl[11:0];
  assign nl_Accum2_acc_92_psp_sva_1 = Accum2_acc_1428_nl + Accum2_acc_1427_nl;
  assign Accum2_acc_92_psp_sva_1 = nl_Accum2_acc_92_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 = (Accum2_acc_93_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[789:785]));
  assign Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1109:1105]));
  assign Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1429:1425]));
  assign Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1749:1745]));
  assign Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1440_nl = conv_s2s_11_12(Product1_3_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1440_nl = nl_Accum2_acc_1440_nl[11:0];
  assign nl_Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4629:4625]));
  assign Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1429_nl = Product1_15_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[149:145]);
  assign Accum2_acc_1429_nl = nl_Accum2_acc_1429_nl[10:0];
  assign nl_Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4949:4945]));
  assign Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[149:145]));
  assign Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[469:465]));
  assign Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1443_nl = Accum2_acc_1440_nl + conv_s2s_11_12(Accum2_acc_1429_nl)
      + conv_s2s_11_12(Product1_16_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1443_nl = nl_Accum2_acc_1443_nl[11:0];
  assign nl_Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3349:3345]));
  assign Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3669:3665]));
  assign Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3989:3985]));
  assign Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4309:4305]));
  assign Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1438_nl = conv_s2s_11_12(Product1_11_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1438_nl = nl_Accum2_acc_1438_nl[11:0];
  assign nl_Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2069:2065]));
  assign Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2389:2385]));
  assign Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2709:2705]));
  assign Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3029:3025]));
  assign Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1442_nl = Accum2_acc_1438_nl + conv_s2s_11_12(Product1_7_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_30_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1442_nl = nl_Accum2_acc_1442_nl[11:0];
  assign nl_Accum2_acc_93_psp_sva_1 = Accum2_acc_1443_nl + Accum2_acc_1442_nl;
  assign Accum2_acc_93_psp_sva_1 = nl_Accum2_acc_93_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 = (Accum2_acc_94_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[794:790]));
  assign Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1114:1110]));
  assign Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1434:1430]));
  assign Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1754:1750]));
  assign Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1455_nl = conv_s2s_11_12(Product1_3_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1455_nl = nl_Accum2_acc_1455_nl[11:0];
  assign nl_Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4634:4630]));
  assign Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1444_nl = Product1_15_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[154:150]);
  assign Accum2_acc_1444_nl = nl_Accum2_acc_1444_nl[10:0];
  assign nl_Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4954:4950]));
  assign Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[154:150]));
  assign Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[474:470]));
  assign Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1458_nl = Accum2_acc_1455_nl + conv_s2s_11_12(Accum2_acc_1444_nl)
      + conv_s2s_11_12(Product1_16_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1458_nl = nl_Accum2_acc_1458_nl[11:0];
  assign nl_Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3354:3350]));
  assign Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3674:3670]));
  assign Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3994:3990]));
  assign Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4314:4310]));
  assign Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1453_nl = conv_s2s_11_12(Product1_11_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1453_nl = nl_Accum2_acc_1453_nl[11:0];
  assign nl_Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2074:2070]));
  assign Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2394:2390]));
  assign Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2714:2710]));
  assign Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3034:3030]));
  assign Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1457_nl = Accum2_acc_1453_nl + conv_s2s_11_12(Product1_7_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_31_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1457_nl = nl_Accum2_acc_1457_nl[11:0];
  assign nl_Accum2_acc_94_psp_sva_1 = Accum2_acc_1458_nl + Accum2_acc_1457_nl;
  assign Accum2_acc_94_psp_sva_1 = nl_Accum2_acc_94_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 = (Accum2_acc_95_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[799:795]));
  assign Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1119:1115]));
  assign Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1439:1435]));
  assign Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1759:1755]));
  assign Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1470_nl = conv_s2s_11_12(Product1_3_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1470_nl = nl_Accum2_acc_1470_nl[11:0];
  assign nl_Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4639:4635]));
  assign Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1459_nl = Product1_15_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[159:155]);
  assign Accum2_acc_1459_nl = nl_Accum2_acc_1459_nl[10:0];
  assign nl_Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4959:4955]));
  assign Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[159:155]));
  assign Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[479:475]));
  assign Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1473_nl = Accum2_acc_1470_nl + conv_s2s_11_12(Accum2_acc_1459_nl)
      + conv_s2s_11_12(Product1_16_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1473_nl = nl_Accum2_acc_1473_nl[11:0];
  assign nl_Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3359:3355]));
  assign Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3679:3675]));
  assign Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[3999:3995]));
  assign Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4319:4315]));
  assign Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1468_nl = conv_s2s_11_12(Product1_11_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1468_nl = nl_Accum2_acc_1468_nl[11:0];
  assign nl_Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2079:2075]));
  assign Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2399:2395]));
  assign Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2719:2715]));
  assign Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3039:3035]));
  assign Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1472_nl = Accum2_acc_1468_nl + conv_s2s_11_12(Product1_7_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_32_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1472_nl = nl_Accum2_acc_1472_nl[11:0];
  assign nl_Accum2_acc_95_psp_sva_1 = Accum2_acc_1473_nl + Accum2_acc_1472_nl;
  assign Accum2_acc_95_psp_sva_1 = nl_Accum2_acc_95_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 = (Accum2_acc_96_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[804:800]));
  assign Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1124:1120]));
  assign Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1444:1440]));
  assign Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1764:1760]));
  assign Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1485_nl = conv_s2s_11_12(Product1_3_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1485_nl = nl_Accum2_acc_1485_nl[11:0];
  assign nl_Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4644:4640]));
  assign Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1474_nl = Product1_15_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[164:160]);
  assign Accum2_acc_1474_nl = nl_Accum2_acc_1474_nl[10:0];
  assign nl_Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4964:4960]));
  assign Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[164:160]));
  assign Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[484:480]));
  assign Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1488_nl = Accum2_acc_1485_nl + conv_s2s_11_12(Accum2_acc_1474_nl)
      + conv_s2s_11_12(Product1_16_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1488_nl = nl_Accum2_acc_1488_nl[11:0];
  assign nl_Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3364:3360]));
  assign Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3684:3680]));
  assign Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4004:4000]));
  assign Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4324:4320]));
  assign Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1483_nl = conv_s2s_11_12(Product1_11_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1483_nl = nl_Accum2_acc_1483_nl[11:0];
  assign nl_Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2084:2080]));
  assign Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2404:2400]));
  assign Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2724:2720]));
  assign Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3044:3040]));
  assign Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1487_nl = Accum2_acc_1483_nl + conv_s2s_11_12(Product1_7_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_33_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1487_nl = nl_Accum2_acc_1487_nl[11:0];
  assign nl_Accum2_acc_96_psp_sva_1 = Accum2_acc_1488_nl + Accum2_acc_1487_nl;
  assign Accum2_acc_96_psp_sva_1 = nl_Accum2_acc_96_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 = (Accum2_acc_97_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[809:805]));
  assign Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1129:1125]));
  assign Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1449:1445]));
  assign Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1769:1765]));
  assign Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1500_nl = conv_s2s_11_12(Product1_3_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1500_nl = nl_Accum2_acc_1500_nl[11:0];
  assign nl_Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4649:4645]));
  assign Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1489_nl = Product1_15_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[169:165]);
  assign Accum2_acc_1489_nl = nl_Accum2_acc_1489_nl[10:0];
  assign nl_Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4969:4965]));
  assign Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[169:165]));
  assign Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[489:485]));
  assign Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1503_nl = Accum2_acc_1500_nl + conv_s2s_11_12(Accum2_acc_1489_nl)
      + conv_s2s_11_12(Product1_16_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1503_nl = nl_Accum2_acc_1503_nl[11:0];
  assign nl_Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3369:3365]));
  assign Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3689:3685]));
  assign Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4009:4005]));
  assign Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4329:4325]));
  assign Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1498_nl = conv_s2s_11_12(Product1_11_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1498_nl = nl_Accum2_acc_1498_nl[11:0];
  assign nl_Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2089:2085]));
  assign Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2409:2405]));
  assign Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2729:2725]));
  assign Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3049:3045]));
  assign Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1502_nl = Accum2_acc_1498_nl + conv_s2s_11_12(Product1_7_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_34_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1502_nl = nl_Accum2_acc_1502_nl[11:0];
  assign nl_Accum2_acc_97_psp_sva_1 = Accum2_acc_1503_nl + Accum2_acc_1502_nl;
  assign Accum2_acc_97_psp_sva_1 = nl_Accum2_acc_97_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 = (Accum2_acc_98_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[814:810]));
  assign Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1134:1130]));
  assign Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1454:1450]));
  assign Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1774:1770]));
  assign Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1515_nl = conv_s2s_11_12(Product1_3_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1515_nl = nl_Accum2_acc_1515_nl[11:0];
  assign nl_Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4654:4650]));
  assign Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1504_nl = Product1_15_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[174:170]);
  assign Accum2_acc_1504_nl = nl_Accum2_acc_1504_nl[10:0];
  assign nl_Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4974:4970]));
  assign Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[174:170]));
  assign Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[494:490]));
  assign Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1518_nl = Accum2_acc_1515_nl + conv_s2s_11_12(Accum2_acc_1504_nl)
      + conv_s2s_11_12(Product1_16_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1518_nl = nl_Accum2_acc_1518_nl[11:0];
  assign nl_Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3374:3370]));
  assign Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3694:3690]));
  assign Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4014:4010]));
  assign Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4334:4330]));
  assign Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1513_nl = conv_s2s_11_12(Product1_11_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1513_nl = nl_Accum2_acc_1513_nl[11:0];
  assign nl_Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2094:2090]));
  assign Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2414:2410]));
  assign Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2734:2730]));
  assign Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3054:3050]));
  assign Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1517_nl = Accum2_acc_1513_nl + conv_s2s_11_12(Product1_7_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_35_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1517_nl = nl_Accum2_acc_1517_nl[11:0];
  assign nl_Accum2_acc_98_psp_sva_1 = Accum2_acc_1518_nl + Accum2_acc_1517_nl;
  assign Accum2_acc_98_psp_sva_1 = nl_Accum2_acc_98_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 = (Accum2_acc_99_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[819:815]));
  assign Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1139:1135]));
  assign Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1459:1455]));
  assign Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1779:1775]));
  assign Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1530_nl = conv_s2s_11_12(Product1_3_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1530_nl = nl_Accum2_acc_1530_nl[11:0];
  assign nl_Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4659:4655]));
  assign Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1519_nl = Product1_15_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[179:175]);
  assign Accum2_acc_1519_nl = nl_Accum2_acc_1519_nl[10:0];
  assign nl_Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4979:4975]));
  assign Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[179:175]));
  assign Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[499:495]));
  assign Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1533_nl = Accum2_acc_1530_nl + conv_s2s_11_12(Accum2_acc_1519_nl)
      + conv_s2s_11_12(Product1_16_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1533_nl = nl_Accum2_acc_1533_nl[11:0];
  assign nl_Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3379:3375]));
  assign Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3699:3695]));
  assign Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4019:4015]));
  assign Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4339:4335]));
  assign Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1528_nl = conv_s2s_11_12(Product1_11_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1528_nl = nl_Accum2_acc_1528_nl[11:0];
  assign nl_Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2099:2095]));
  assign Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2419:2415]));
  assign Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2739:2735]));
  assign Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3059:3055]));
  assign Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1532_nl = Accum2_acc_1528_nl + conv_s2s_11_12(Product1_7_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_36_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1532_nl = nl_Accum2_acc_1532_nl[11:0];
  assign nl_Accum2_acc_99_psp_sva_1 = Accum2_acc_1533_nl + Accum2_acc_1532_nl;
  assign Accum2_acc_99_psp_sva_1 = nl_Accum2_acc_99_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 = (Accum2_acc_100_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[824:820]));
  assign Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1144:1140]));
  assign Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1464:1460]));
  assign Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1784:1780]));
  assign Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1545_nl = conv_s2s_11_12(Product1_3_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1545_nl = nl_Accum2_acc_1545_nl[11:0];
  assign nl_Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4664:4660]));
  assign Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1534_nl = Product1_15_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[184:180]);
  assign Accum2_acc_1534_nl = nl_Accum2_acc_1534_nl[10:0];
  assign nl_Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4984:4980]));
  assign Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[184:180]));
  assign Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[504:500]));
  assign Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1548_nl = Accum2_acc_1545_nl + conv_s2s_11_12(Accum2_acc_1534_nl)
      + conv_s2s_11_12(Product1_16_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1548_nl = nl_Accum2_acc_1548_nl[11:0];
  assign nl_Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3384:3380]));
  assign Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3704:3700]));
  assign Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4024:4020]));
  assign Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4344:4340]));
  assign Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1543_nl = conv_s2s_11_12(Product1_11_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1543_nl = nl_Accum2_acc_1543_nl[11:0];
  assign nl_Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2104:2100]));
  assign Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2424:2420]));
  assign Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2744:2740]));
  assign Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3064:3060]));
  assign Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1547_nl = Accum2_acc_1543_nl + conv_s2s_11_12(Product1_7_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_37_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1547_nl = nl_Accum2_acc_1547_nl[11:0];
  assign nl_Accum2_acc_100_psp_sva_1 = Accum2_acc_1548_nl + Accum2_acc_1547_nl;
  assign Accum2_acc_100_psp_sva_1 = nl_Accum2_acc_100_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 = (Accum2_acc_101_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[829:825]));
  assign Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1149:1145]));
  assign Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1469:1465]));
  assign Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1789:1785]));
  assign Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1560_nl = conv_s2s_11_12(Product1_3_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1560_nl = nl_Accum2_acc_1560_nl[11:0];
  assign nl_Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4669:4665]));
  assign Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1549_nl = Product1_15_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[189:185]);
  assign Accum2_acc_1549_nl = nl_Accum2_acc_1549_nl[10:0];
  assign nl_Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4989:4985]));
  assign Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[189:185]));
  assign Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[509:505]));
  assign Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1563_nl = Accum2_acc_1560_nl + conv_s2s_11_12(Accum2_acc_1549_nl)
      + conv_s2s_11_12(Product1_16_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1563_nl = nl_Accum2_acc_1563_nl[11:0];
  assign nl_Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3389:3385]));
  assign Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3709:3705]));
  assign Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4029:4025]));
  assign Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4349:4345]));
  assign Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1558_nl = conv_s2s_11_12(Product1_11_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1558_nl = nl_Accum2_acc_1558_nl[11:0];
  assign nl_Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2109:2105]));
  assign Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2429:2425]));
  assign Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2749:2745]));
  assign Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3069:3065]));
  assign Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1562_nl = Accum2_acc_1558_nl + conv_s2s_11_12(Product1_7_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_38_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1562_nl = nl_Accum2_acc_1562_nl[11:0];
  assign nl_Accum2_acc_101_psp_sva_1 = Accum2_acc_1563_nl + Accum2_acc_1562_nl;
  assign Accum2_acc_101_psp_sva_1 = nl_Accum2_acc_101_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 = (Accum2_acc_102_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[834:830]));
  assign Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1154:1150]));
  assign Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1474:1470]));
  assign Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1794:1790]));
  assign Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1575_nl = conv_s2s_11_12(Product1_3_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1575_nl = nl_Accum2_acc_1575_nl[11:0];
  assign nl_Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4674:4670]));
  assign Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1564_nl = Product1_15_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[194:190]);
  assign Accum2_acc_1564_nl = nl_Accum2_acc_1564_nl[10:0];
  assign nl_Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4994:4990]));
  assign Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[194:190]));
  assign Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[514:510]));
  assign Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1578_nl = Accum2_acc_1575_nl + conv_s2s_11_12(Accum2_acc_1564_nl)
      + conv_s2s_11_12(Product1_16_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1578_nl = nl_Accum2_acc_1578_nl[11:0];
  assign nl_Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3394:3390]));
  assign Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3714:3710]));
  assign Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4034:4030]));
  assign Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4354:4350]));
  assign Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1573_nl = conv_s2s_11_12(Product1_11_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1573_nl = nl_Accum2_acc_1573_nl[11:0];
  assign nl_Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2114:2110]));
  assign Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2434:2430]));
  assign Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2754:2750]));
  assign Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3074:3070]));
  assign Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1577_nl = Accum2_acc_1573_nl + conv_s2s_11_12(Product1_7_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_39_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1577_nl = nl_Accum2_acc_1577_nl[11:0];
  assign nl_Accum2_acc_102_psp_sva_1 = Accum2_acc_1578_nl + Accum2_acc_1577_nl;
  assign Accum2_acc_102_psp_sva_1 = nl_Accum2_acc_102_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 = (Accum2_acc_103_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[839:835]));
  assign Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1159:1155]));
  assign Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1479:1475]));
  assign Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1799:1795]));
  assign Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1590_nl = conv_s2s_11_12(Product1_3_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1590_nl = nl_Accum2_acc_1590_nl[11:0];
  assign nl_Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4679:4675]));
  assign Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1579_nl = Product1_15_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[199:195]);
  assign Accum2_acc_1579_nl = nl_Accum2_acc_1579_nl[10:0];
  assign nl_Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[4999:4995]));
  assign Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[199:195]));
  assign Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[519:515]));
  assign Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1593_nl = Accum2_acc_1590_nl + conv_s2s_11_12(Accum2_acc_1579_nl)
      + conv_s2s_11_12(Product1_16_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1593_nl = nl_Accum2_acc_1593_nl[11:0];
  assign nl_Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3399:3395]));
  assign Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3719:3715]));
  assign Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4039:4035]));
  assign Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4359:4355]));
  assign Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1588_nl = conv_s2s_11_12(Product1_11_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1588_nl = nl_Accum2_acc_1588_nl[11:0];
  assign nl_Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2119:2115]));
  assign Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2439:2435]));
  assign Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2759:2755]));
  assign Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3079:3075]));
  assign Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1592_nl = Accum2_acc_1588_nl + conv_s2s_11_12(Product1_7_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_40_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1592_nl = nl_Accum2_acc_1592_nl[11:0];
  assign nl_Accum2_acc_103_psp_sva_1 = Accum2_acc_1593_nl + Accum2_acc_1592_nl;
  assign Accum2_acc_103_psp_sva_1 = nl_Accum2_acc_103_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 = (Accum2_acc_104_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[844:840]));
  assign Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1164:1160]));
  assign Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1484:1480]));
  assign Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1804:1800]));
  assign Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1605_nl = conv_s2s_11_12(Product1_3_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1605_nl = nl_Accum2_acc_1605_nl[11:0];
  assign nl_Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4684:4680]));
  assign Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1594_nl = Product1_15_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[204:200]);
  assign Accum2_acc_1594_nl = nl_Accum2_acc_1594_nl[10:0];
  assign nl_Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5004:5000]));
  assign Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[204:200]));
  assign Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[524:520]));
  assign Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1608_nl = Accum2_acc_1605_nl + conv_s2s_11_12(Accum2_acc_1594_nl)
      + conv_s2s_11_12(Product1_16_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1608_nl = nl_Accum2_acc_1608_nl[11:0];
  assign nl_Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3404:3400]));
  assign Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3724:3720]));
  assign Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4044:4040]));
  assign Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4364:4360]));
  assign Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1603_nl = conv_s2s_11_12(Product1_11_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1603_nl = nl_Accum2_acc_1603_nl[11:0];
  assign nl_Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2124:2120]));
  assign Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2444:2440]));
  assign Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2764:2760]));
  assign Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3084:3080]));
  assign Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1607_nl = Accum2_acc_1603_nl + conv_s2s_11_12(Product1_7_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_41_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1607_nl = nl_Accum2_acc_1607_nl[11:0];
  assign nl_Accum2_acc_104_psp_sva_1 = Accum2_acc_1608_nl + Accum2_acc_1607_nl;
  assign Accum2_acc_104_psp_sva_1 = nl_Accum2_acc_104_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 = (Accum2_acc_105_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[849:845]));
  assign Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1169:1165]));
  assign Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1489:1485]));
  assign Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1809:1805]));
  assign Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1620_nl = conv_s2s_11_12(Product1_3_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1620_nl = nl_Accum2_acc_1620_nl[11:0];
  assign nl_Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4689:4685]));
  assign Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1609_nl = Product1_15_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[209:205]);
  assign Accum2_acc_1609_nl = nl_Accum2_acc_1609_nl[10:0];
  assign nl_Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5009:5005]));
  assign Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[209:205]));
  assign Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[529:525]));
  assign Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1623_nl = Accum2_acc_1620_nl + conv_s2s_11_12(Accum2_acc_1609_nl)
      + conv_s2s_11_12(Product1_16_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1623_nl = nl_Accum2_acc_1623_nl[11:0];
  assign nl_Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3409:3405]));
  assign Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3729:3725]));
  assign Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4049:4045]));
  assign Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4369:4365]));
  assign Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1618_nl = conv_s2s_11_12(Product1_11_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1618_nl = nl_Accum2_acc_1618_nl[11:0];
  assign nl_Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2129:2125]));
  assign Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2449:2445]));
  assign Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2769:2765]));
  assign Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3089:3085]));
  assign Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1622_nl = Accum2_acc_1618_nl + conv_s2s_11_12(Product1_7_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_42_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1622_nl = nl_Accum2_acc_1622_nl[11:0];
  assign nl_Accum2_acc_105_psp_sva_1 = Accum2_acc_1623_nl + Accum2_acc_1622_nl;
  assign Accum2_acc_105_psp_sva_1 = nl_Accum2_acc_105_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 = (Accum2_acc_106_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[854:850]));
  assign Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1174:1170]));
  assign Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1494:1490]));
  assign Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1814:1810]));
  assign Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1635_nl = conv_s2s_11_12(Product1_3_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1635_nl = nl_Accum2_acc_1635_nl[11:0];
  assign nl_Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4694:4690]));
  assign Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1624_nl = Product1_15_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[214:210]);
  assign Accum2_acc_1624_nl = nl_Accum2_acc_1624_nl[10:0];
  assign nl_Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5014:5010]));
  assign Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[214:210]));
  assign Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[534:530]));
  assign Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1638_nl = Accum2_acc_1635_nl + conv_s2s_11_12(Accum2_acc_1624_nl)
      + conv_s2s_11_12(Product1_16_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1638_nl = nl_Accum2_acc_1638_nl[11:0];
  assign nl_Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3414:3410]));
  assign Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3734:3730]));
  assign Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4054:4050]));
  assign Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4374:4370]));
  assign Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1633_nl = conv_s2s_11_12(Product1_11_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1633_nl = nl_Accum2_acc_1633_nl[11:0];
  assign nl_Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2134:2130]));
  assign Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2454:2450]));
  assign Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2774:2770]));
  assign Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3094:3090]));
  assign Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1637_nl = Accum2_acc_1633_nl + conv_s2s_11_12(Product1_7_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_43_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1637_nl = nl_Accum2_acc_1637_nl[11:0];
  assign nl_Accum2_acc_106_psp_sva_1 = Accum2_acc_1638_nl + Accum2_acc_1637_nl;
  assign Accum2_acc_106_psp_sva_1 = nl_Accum2_acc_106_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 = (Accum2_acc_107_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[859:855]));
  assign Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1179:1175]));
  assign Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1499:1495]));
  assign Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1819:1815]));
  assign Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1650_nl = conv_s2s_11_12(Product1_3_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1650_nl = nl_Accum2_acc_1650_nl[11:0];
  assign nl_Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4699:4695]));
  assign Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1639_nl = Product1_15_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[219:215]);
  assign Accum2_acc_1639_nl = nl_Accum2_acc_1639_nl[10:0];
  assign nl_Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5019:5015]));
  assign Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[219:215]));
  assign Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[539:535]));
  assign Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1653_nl = Accum2_acc_1650_nl + conv_s2s_11_12(Accum2_acc_1639_nl)
      + conv_s2s_11_12(Product1_16_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1653_nl = nl_Accum2_acc_1653_nl[11:0];
  assign nl_Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3419:3415]));
  assign Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3739:3735]));
  assign Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4059:4055]));
  assign Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4379:4375]));
  assign Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1648_nl = conv_s2s_11_12(Product1_11_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1648_nl = nl_Accum2_acc_1648_nl[11:0];
  assign nl_Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2139:2135]));
  assign Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2459:2455]));
  assign Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2779:2775]));
  assign Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3099:3095]));
  assign Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1652_nl = Accum2_acc_1648_nl + conv_s2s_11_12(Product1_7_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_44_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1652_nl = nl_Accum2_acc_1652_nl[11:0];
  assign nl_Accum2_acc_107_psp_sva_1 = Accum2_acc_1653_nl + Accum2_acc_1652_nl;
  assign Accum2_acc_107_psp_sva_1 = nl_Accum2_acc_107_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 = (Accum2_acc_108_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[864:860]));
  assign Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1184:1180]));
  assign Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1504:1500]));
  assign Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1824:1820]));
  assign Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1665_nl = conv_s2s_11_12(Product1_3_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1665_nl = nl_Accum2_acc_1665_nl[11:0];
  assign nl_Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4704:4700]));
  assign Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1654_nl = Product1_15_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[224:220]);
  assign Accum2_acc_1654_nl = nl_Accum2_acc_1654_nl[10:0];
  assign nl_Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5024:5020]));
  assign Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[224:220]));
  assign Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[544:540]));
  assign Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1668_nl = Accum2_acc_1665_nl + conv_s2s_11_12(Accum2_acc_1654_nl)
      + conv_s2s_11_12(Product1_16_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1668_nl = nl_Accum2_acc_1668_nl[11:0];
  assign nl_Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3424:3420]));
  assign Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3744:3740]));
  assign Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4064:4060]));
  assign Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4384:4380]));
  assign Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1663_nl = conv_s2s_11_12(Product1_11_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1663_nl = nl_Accum2_acc_1663_nl[11:0];
  assign nl_Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2144:2140]));
  assign Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2464:2460]));
  assign Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2784:2780]));
  assign Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3104:3100]));
  assign Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1667_nl = Accum2_acc_1663_nl + conv_s2s_11_12(Product1_7_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_45_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1667_nl = nl_Accum2_acc_1667_nl[11:0];
  assign nl_Accum2_acc_108_psp_sva_1 = Accum2_acc_1668_nl + Accum2_acc_1667_nl;
  assign Accum2_acc_108_psp_sva_1 = nl_Accum2_acc_108_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 = (Accum2_acc_109_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[869:865]));
  assign Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1189:1185]));
  assign Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1509:1505]));
  assign Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1829:1825]));
  assign Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1680_nl = conv_s2s_11_12(Product1_3_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1680_nl = nl_Accum2_acc_1680_nl[11:0];
  assign nl_Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4709:4705]));
  assign Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1669_nl = Product1_15_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[229:225]);
  assign Accum2_acc_1669_nl = nl_Accum2_acc_1669_nl[10:0];
  assign nl_Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5029:5025]));
  assign Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[229:225]));
  assign Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[549:545]));
  assign Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1683_nl = Accum2_acc_1680_nl + conv_s2s_11_12(Accum2_acc_1669_nl)
      + conv_s2s_11_12(Product1_16_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1683_nl = nl_Accum2_acc_1683_nl[11:0];
  assign nl_Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3429:3425]));
  assign Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3749:3745]));
  assign Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4069:4065]));
  assign Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4389:4385]));
  assign Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1678_nl = conv_s2s_11_12(Product1_11_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1678_nl = nl_Accum2_acc_1678_nl[11:0];
  assign nl_Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2149:2145]));
  assign Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2469:2465]));
  assign Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2789:2785]));
  assign Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3109:3105]));
  assign Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1682_nl = Accum2_acc_1678_nl + conv_s2s_11_12(Product1_7_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_46_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1682_nl = nl_Accum2_acc_1682_nl[11:0];
  assign nl_Accum2_acc_109_psp_sva_1 = Accum2_acc_1683_nl + Accum2_acc_1682_nl;
  assign Accum2_acc_109_psp_sva_1 = nl_Accum2_acc_109_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 = (Accum2_acc_110_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[874:870]));
  assign Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1194:1190]));
  assign Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1514:1510]));
  assign Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1834:1830]));
  assign Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1695_nl = conv_s2s_11_12(Product1_3_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1695_nl = nl_Accum2_acc_1695_nl[11:0];
  assign nl_Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4714:4710]));
  assign Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1684_nl = Product1_15_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[234:230]);
  assign Accum2_acc_1684_nl = nl_Accum2_acc_1684_nl[10:0];
  assign nl_Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5034:5030]));
  assign Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[234:230]));
  assign Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[554:550]));
  assign Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1698_nl = Accum2_acc_1695_nl + conv_s2s_11_12(Accum2_acc_1684_nl)
      + conv_s2s_11_12(Product1_16_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1698_nl = nl_Accum2_acc_1698_nl[11:0];
  assign nl_Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3434:3430]));
  assign Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3754:3750]));
  assign Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4074:4070]));
  assign Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4394:4390]));
  assign Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1693_nl = conv_s2s_11_12(Product1_11_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1693_nl = nl_Accum2_acc_1693_nl[11:0];
  assign nl_Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2154:2150]));
  assign Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2474:2470]));
  assign Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2794:2790]));
  assign Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3114:3110]));
  assign Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1697_nl = Accum2_acc_1693_nl + conv_s2s_11_12(Product1_7_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_47_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1697_nl = nl_Accum2_acc_1697_nl[11:0];
  assign nl_Accum2_acc_110_psp_sva_1 = Accum2_acc_1698_nl + Accum2_acc_1697_nl;
  assign Accum2_acc_110_psp_sva_1 = nl_Accum2_acc_110_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 = (Accum2_acc_111_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[879:875]));
  assign Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1199:1195]));
  assign Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1519:1515]));
  assign Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1839:1835]));
  assign Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1710_nl = conv_s2s_11_12(Product1_3_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1710_nl = nl_Accum2_acc_1710_nl[11:0];
  assign nl_Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4719:4715]));
  assign Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1699_nl = Product1_15_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[239:235]);
  assign Accum2_acc_1699_nl = nl_Accum2_acc_1699_nl[10:0];
  assign nl_Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5039:5035]));
  assign Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[239:235]));
  assign Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[559:555]));
  assign Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1713_nl = Accum2_acc_1710_nl + conv_s2s_11_12(Accum2_acc_1699_nl)
      + conv_s2s_11_12(Product1_16_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1713_nl = nl_Accum2_acc_1713_nl[11:0];
  assign nl_Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3439:3435]));
  assign Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3759:3755]));
  assign Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4079:4075]));
  assign Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4399:4395]));
  assign Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1708_nl = conv_s2s_11_12(Product1_11_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1708_nl = nl_Accum2_acc_1708_nl[11:0];
  assign nl_Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2159:2155]));
  assign Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2479:2475]));
  assign Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2799:2795]));
  assign Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3119:3115]));
  assign Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1712_nl = Accum2_acc_1708_nl + conv_s2s_11_12(Product1_7_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_48_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1712_nl = nl_Accum2_acc_1712_nl[11:0];
  assign nl_Accum2_acc_111_psp_sva_1 = Accum2_acc_1713_nl + Accum2_acc_1712_nl;
  assign Accum2_acc_111_psp_sva_1 = nl_Accum2_acc_111_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 = (Accum2_acc_112_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[884:880]));
  assign Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1204:1200]));
  assign Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1524:1520]));
  assign Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1844:1840]));
  assign Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1725_nl = conv_s2s_11_12(Product1_3_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1725_nl = nl_Accum2_acc_1725_nl[11:0];
  assign nl_Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4724:4720]));
  assign Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1714_nl = Product1_15_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[244:240]);
  assign Accum2_acc_1714_nl = nl_Accum2_acc_1714_nl[10:0];
  assign nl_Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5044:5040]));
  assign Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[244:240]));
  assign Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[564:560]));
  assign Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1728_nl = Accum2_acc_1725_nl + conv_s2s_11_12(Accum2_acc_1714_nl)
      + conv_s2s_11_12(Product1_16_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1728_nl = nl_Accum2_acc_1728_nl[11:0];
  assign nl_Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3444:3440]));
  assign Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3764:3760]));
  assign Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4084:4080]));
  assign Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4404:4400]));
  assign Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1723_nl = conv_s2s_11_12(Product1_11_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1723_nl = nl_Accum2_acc_1723_nl[11:0];
  assign nl_Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2164:2160]));
  assign Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2484:2480]));
  assign Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2804:2800]));
  assign Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3124:3120]));
  assign Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1727_nl = Accum2_acc_1723_nl + conv_s2s_11_12(Product1_7_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_49_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1727_nl = nl_Accum2_acc_1727_nl[11:0];
  assign nl_Accum2_acc_112_psp_sva_1 = Accum2_acc_1728_nl + Accum2_acc_1727_nl;
  assign Accum2_acc_112_psp_sva_1 = nl_Accum2_acc_112_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 = (Accum2_acc_113_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[889:885]));
  assign Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1209:1205]));
  assign Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1529:1525]));
  assign Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1849:1845]));
  assign Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1740_nl = conv_s2s_11_12(Product1_3_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1740_nl = nl_Accum2_acc_1740_nl[11:0];
  assign nl_Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4729:4725]));
  assign Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1729_nl = Product1_15_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[249:245]);
  assign Accum2_acc_1729_nl = nl_Accum2_acc_1729_nl[10:0];
  assign nl_Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5049:5045]));
  assign Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[249:245]));
  assign Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[569:565]));
  assign Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1743_nl = Accum2_acc_1740_nl + conv_s2s_11_12(Accum2_acc_1729_nl)
      + conv_s2s_11_12(Product1_16_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1743_nl = nl_Accum2_acc_1743_nl[11:0];
  assign nl_Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3449:3445]));
  assign Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3769:3765]));
  assign Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4089:4085]));
  assign Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4409:4405]));
  assign Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1738_nl = conv_s2s_11_12(Product1_11_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1738_nl = nl_Accum2_acc_1738_nl[11:0];
  assign nl_Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2169:2165]));
  assign Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2489:2485]));
  assign Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2809:2805]));
  assign Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3129:3125]));
  assign Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1742_nl = Accum2_acc_1738_nl + conv_s2s_11_12(Product1_7_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_50_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1742_nl = nl_Accum2_acc_1742_nl[11:0];
  assign nl_Accum2_acc_113_psp_sva_1 = Accum2_acc_1743_nl + Accum2_acc_1742_nl;
  assign Accum2_acc_113_psp_sva_1 = nl_Accum2_acc_113_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 = (Accum2_acc_114_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[894:890]));
  assign Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1214:1210]));
  assign Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1534:1530]));
  assign Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1854:1850]));
  assign Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1755_nl = conv_s2s_11_12(Product1_3_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1755_nl = nl_Accum2_acc_1755_nl[11:0];
  assign nl_Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4734:4730]));
  assign Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1744_nl = Product1_15_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[254:250]);
  assign Accum2_acc_1744_nl = nl_Accum2_acc_1744_nl[10:0];
  assign nl_Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5054:5050]));
  assign Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[254:250]));
  assign Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[574:570]));
  assign Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1758_nl = Accum2_acc_1755_nl + conv_s2s_11_12(Accum2_acc_1744_nl)
      + conv_s2s_11_12(Product1_16_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1758_nl = nl_Accum2_acc_1758_nl[11:0];
  assign nl_Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3454:3450]));
  assign Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3774:3770]));
  assign Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4094:4090]));
  assign Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4414:4410]));
  assign Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1753_nl = conv_s2s_11_12(Product1_11_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1753_nl = nl_Accum2_acc_1753_nl[11:0];
  assign nl_Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2174:2170]));
  assign Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2494:2490]));
  assign Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2814:2810]));
  assign Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3134:3130]));
  assign Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1757_nl = Accum2_acc_1753_nl + conv_s2s_11_12(Product1_7_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_51_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1757_nl = nl_Accum2_acc_1757_nl[11:0];
  assign nl_Accum2_acc_114_psp_sva_1 = Accum2_acc_1758_nl + Accum2_acc_1757_nl;
  assign Accum2_acc_114_psp_sva_1 = nl_Accum2_acc_114_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 = (Accum2_acc_115_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[899:895]));
  assign Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1219:1215]));
  assign Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1539:1535]));
  assign Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1859:1855]));
  assign Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1770_nl = conv_s2s_11_12(Product1_3_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1770_nl = nl_Accum2_acc_1770_nl[11:0];
  assign nl_Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4739:4735]));
  assign Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1759_nl = Product1_15_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[259:255]);
  assign Accum2_acc_1759_nl = nl_Accum2_acc_1759_nl[10:0];
  assign nl_Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5059:5055]));
  assign Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[259:255]));
  assign Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[579:575]));
  assign Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1773_nl = Accum2_acc_1770_nl + conv_s2s_11_12(Accum2_acc_1759_nl)
      + conv_s2s_11_12(Product1_16_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1773_nl = nl_Accum2_acc_1773_nl[11:0];
  assign nl_Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3459:3455]));
  assign Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3779:3775]));
  assign Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4099:4095]));
  assign Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4419:4415]));
  assign Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1768_nl = conv_s2s_11_12(Product1_11_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1768_nl = nl_Accum2_acc_1768_nl[11:0];
  assign nl_Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2179:2175]));
  assign Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2499:2495]));
  assign Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2819:2815]));
  assign Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3139:3135]));
  assign Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1772_nl = Accum2_acc_1768_nl + conv_s2s_11_12(Product1_7_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_52_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1772_nl = nl_Accum2_acc_1772_nl[11:0];
  assign nl_Accum2_acc_115_psp_sva_1 = Accum2_acc_1773_nl + Accum2_acc_1772_nl;
  assign Accum2_acc_115_psp_sva_1 = nl_Accum2_acc_115_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 = (Accum2_acc_116_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[904:900]));
  assign Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1224:1220]));
  assign Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1544:1540]));
  assign Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1864:1860]));
  assign Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1785_nl = conv_s2s_11_12(Product1_3_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1785_nl = nl_Accum2_acc_1785_nl[11:0];
  assign nl_Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4744:4740]));
  assign Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1774_nl = Product1_15_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[264:260]);
  assign Accum2_acc_1774_nl = nl_Accum2_acc_1774_nl[10:0];
  assign nl_Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5064:5060]));
  assign Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[264:260]));
  assign Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[584:580]));
  assign Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1788_nl = Accum2_acc_1785_nl + conv_s2s_11_12(Accum2_acc_1774_nl)
      + conv_s2s_11_12(Product1_16_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1788_nl = nl_Accum2_acc_1788_nl[11:0];
  assign nl_Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3464:3460]));
  assign Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3784:3780]));
  assign Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4104:4100]));
  assign Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4424:4420]));
  assign Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1783_nl = conv_s2s_11_12(Product1_11_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1783_nl = nl_Accum2_acc_1783_nl[11:0];
  assign nl_Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2184:2180]));
  assign Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2504:2500]));
  assign Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2824:2820]));
  assign Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3144:3140]));
  assign Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1787_nl = Accum2_acc_1783_nl + conv_s2s_11_12(Product1_7_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_53_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1787_nl = nl_Accum2_acc_1787_nl[11:0];
  assign nl_Accum2_acc_116_psp_sva_1 = Accum2_acc_1788_nl + Accum2_acc_1787_nl;
  assign Accum2_acc_116_psp_sva_1 = nl_Accum2_acc_116_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 = (Accum2_acc_117_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[909:905]));
  assign Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1229:1225]));
  assign Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1549:1545]));
  assign Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1869:1865]));
  assign Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1800_nl = conv_s2s_11_12(Product1_3_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1800_nl = nl_Accum2_acc_1800_nl[11:0];
  assign nl_Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4749:4745]));
  assign Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1789_nl = Product1_15_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[269:265]);
  assign Accum2_acc_1789_nl = nl_Accum2_acc_1789_nl[10:0];
  assign nl_Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5069:5065]));
  assign Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[269:265]));
  assign Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[589:585]));
  assign Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1803_nl = Accum2_acc_1800_nl + conv_s2s_11_12(Accum2_acc_1789_nl)
      + conv_s2s_11_12(Product1_16_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1803_nl = nl_Accum2_acc_1803_nl[11:0];
  assign nl_Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3469:3465]));
  assign Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3789:3785]));
  assign Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4109:4105]));
  assign Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4429:4425]));
  assign Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1798_nl = conv_s2s_11_12(Product1_11_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1798_nl = nl_Accum2_acc_1798_nl[11:0];
  assign nl_Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2189:2185]));
  assign Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2509:2505]));
  assign Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2829:2825]));
  assign Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3149:3145]));
  assign Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1802_nl = Accum2_acc_1798_nl + conv_s2s_11_12(Product1_7_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_54_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1802_nl = nl_Accum2_acc_1802_nl[11:0];
  assign nl_Accum2_acc_117_psp_sva_1 = Accum2_acc_1803_nl + Accum2_acc_1802_nl;
  assign Accum2_acc_117_psp_sva_1 = nl_Accum2_acc_117_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 = (Accum2_acc_118_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[914:910]));
  assign Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1234:1230]));
  assign Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1554:1550]));
  assign Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1874:1870]));
  assign Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1815_nl = conv_s2s_11_12(Product1_3_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1815_nl = nl_Accum2_acc_1815_nl[11:0];
  assign nl_Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4754:4750]));
  assign Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1804_nl = Product1_15_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[274:270]);
  assign Accum2_acc_1804_nl = nl_Accum2_acc_1804_nl[10:0];
  assign nl_Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5074:5070]));
  assign Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[274:270]));
  assign Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[594:590]));
  assign Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1818_nl = Accum2_acc_1815_nl + conv_s2s_11_12(Accum2_acc_1804_nl)
      + conv_s2s_11_12(Product1_16_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1818_nl = nl_Accum2_acc_1818_nl[11:0];
  assign nl_Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3474:3470]));
  assign Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3794:3790]));
  assign Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4114:4110]));
  assign Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4434:4430]));
  assign Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1813_nl = conv_s2s_11_12(Product1_11_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1813_nl = nl_Accum2_acc_1813_nl[11:0];
  assign nl_Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2194:2190]));
  assign Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2514:2510]));
  assign Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2834:2830]));
  assign Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3154:3150]));
  assign Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1817_nl = Accum2_acc_1813_nl + conv_s2s_11_12(Product1_7_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_55_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1817_nl = nl_Accum2_acc_1817_nl[11:0];
  assign nl_Accum2_acc_118_psp_sva_1 = Accum2_acc_1818_nl + Accum2_acc_1817_nl;
  assign Accum2_acc_118_psp_sva_1 = nl_Accum2_acc_118_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 = (Accum2_acc_119_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[919:915]));
  assign Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1239:1235]));
  assign Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1559:1555]));
  assign Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1879:1875]));
  assign Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1830_nl = conv_s2s_11_12(Product1_3_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1830_nl = nl_Accum2_acc_1830_nl[11:0];
  assign nl_Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4759:4755]));
  assign Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1819_nl = Product1_15_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[279:275]);
  assign Accum2_acc_1819_nl = nl_Accum2_acc_1819_nl[10:0];
  assign nl_Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5079:5075]));
  assign Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[279:275]));
  assign Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[599:595]));
  assign Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1833_nl = Accum2_acc_1830_nl + conv_s2s_11_12(Accum2_acc_1819_nl)
      + conv_s2s_11_12(Product1_16_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1833_nl = nl_Accum2_acc_1833_nl[11:0];
  assign nl_Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3479:3475]));
  assign Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3799:3795]));
  assign Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4119:4115]));
  assign Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4439:4435]));
  assign Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1828_nl = conv_s2s_11_12(Product1_11_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1828_nl = nl_Accum2_acc_1828_nl[11:0];
  assign nl_Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2199:2195]));
  assign Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2519:2515]));
  assign Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2839:2835]));
  assign Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3159:3155]));
  assign Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1832_nl = Accum2_acc_1828_nl + conv_s2s_11_12(Product1_7_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_56_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1832_nl = nl_Accum2_acc_1832_nl[11:0];
  assign nl_Accum2_acc_119_psp_sva_1 = Accum2_acc_1833_nl + Accum2_acc_1832_nl;
  assign Accum2_acc_119_psp_sva_1 = nl_Accum2_acc_119_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 = (Accum2_acc_120_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[924:920]));
  assign Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1244:1240]));
  assign Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1564:1560]));
  assign Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1884:1880]));
  assign Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1845_nl = conv_s2s_11_12(Product1_3_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1845_nl = nl_Accum2_acc_1845_nl[11:0];
  assign nl_Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4764:4760]));
  assign Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1834_nl = Product1_15_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[284:280]);
  assign Accum2_acc_1834_nl = nl_Accum2_acc_1834_nl[10:0];
  assign nl_Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5084:5080]));
  assign Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[284:280]));
  assign Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[604:600]));
  assign Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1848_nl = Accum2_acc_1845_nl + conv_s2s_11_12(Accum2_acc_1834_nl)
      + conv_s2s_11_12(Product1_16_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1848_nl = nl_Accum2_acc_1848_nl[11:0];
  assign nl_Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3484:3480]));
  assign Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3804:3800]));
  assign Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4124:4120]));
  assign Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4444:4440]));
  assign Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1843_nl = conv_s2s_11_12(Product1_11_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1843_nl = nl_Accum2_acc_1843_nl[11:0];
  assign nl_Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2204:2200]));
  assign Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2524:2520]));
  assign Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2844:2840]));
  assign Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3164:3160]));
  assign Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1847_nl = Accum2_acc_1843_nl + conv_s2s_11_12(Product1_7_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_57_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1847_nl = nl_Accum2_acc_1847_nl[11:0];
  assign nl_Accum2_acc_120_psp_sva_1 = Accum2_acc_1848_nl + Accum2_acc_1847_nl;
  assign Accum2_acc_120_psp_sva_1 = nl_Accum2_acc_120_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1 = (Accum2_acc_121_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[929:925]));
  assign Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1249:1245]));
  assign Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1569:1565]));
  assign Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1889:1885]));
  assign Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1860_nl = conv_s2s_11_12(Product1_3_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1860_nl = nl_Accum2_acc_1860_nl[11:0];
  assign nl_Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4769:4765]));
  assign Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1849_nl = Product1_15_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[289:285]);
  assign Accum2_acc_1849_nl = nl_Accum2_acc_1849_nl[10:0];
  assign nl_Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5089:5085]));
  assign Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[289:285]));
  assign Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[609:605]));
  assign Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1863_nl = Accum2_acc_1860_nl + conv_s2s_11_12(Accum2_acc_1849_nl)
      + conv_s2s_11_12(Product1_16_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1863_nl = nl_Accum2_acc_1863_nl[11:0];
  assign nl_Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3489:3485]));
  assign Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3809:3805]));
  assign Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4129:4125]));
  assign Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4449:4445]));
  assign Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1858_nl = conv_s2s_11_12(Product1_11_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1858_nl = nl_Accum2_acc_1858_nl[11:0];
  assign nl_Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2209:2205]));
  assign Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2529:2525]));
  assign Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2849:2845]));
  assign Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3169:3165]));
  assign Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1862_nl = Accum2_acc_1858_nl + conv_s2s_11_12(Product1_7_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_58_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1862_nl = nl_Accum2_acc_1862_nl[11:0];
  assign nl_Accum2_acc_121_psp_sva_1 = Accum2_acc_1863_nl + Accum2_acc_1862_nl;
  assign Accum2_acc_121_psp_sva_1 = nl_Accum2_acc_121_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1 = (Accum2_acc_122_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[934:930]));
  assign Product1_3_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1254:1250]));
  assign Product1_4_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1574:1570]));
  assign Product1_5_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1894:1890]));
  assign Product1_6_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1875_nl = conv_s2s_11_12(Product1_3_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1875_nl = nl_Accum2_acc_1875_nl[11:0];
  assign nl_Product1_15_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4774:4770]));
  assign Product1_15_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1864_nl = Product1_15_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[294:290]);
  assign Accum2_acc_1864_nl = nl_Accum2_acc_1864_nl[10:0];
  assign nl_Product1_16_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5094:5090]));
  assign Product1_16_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[294:290]));
  assign Product1_1_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[614:610]));
  assign Product1_2_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1878_nl = Accum2_acc_1875_nl + conv_s2s_11_12(Accum2_acc_1864_nl)
      + conv_s2s_11_12(Product1_16_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1878_nl = nl_Accum2_acc_1878_nl[11:0];
  assign nl_Product1_11_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3494:3490]));
  assign Product1_11_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3814:3810]));
  assign Product1_12_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4134:4130]));
  assign Product1_13_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4454:4450]));
  assign Product1_14_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1873_nl = conv_s2s_11_12(Product1_11_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1873_nl = nl_Accum2_acc_1873_nl[11:0];
  assign nl_Product1_7_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2214:2210]));
  assign Product1_7_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2534:2530]));
  assign Product1_8_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2854:2850]));
  assign Product1_9_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3174:3170]));
  assign Product1_10_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1877_nl = Accum2_acc_1873_nl + conv_s2s_11_12(Product1_7_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_59_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1877_nl = nl_Accum2_acc_1877_nl[11:0];
  assign nl_Accum2_acc_122_psp_sva_1 = Accum2_acc_1878_nl + Accum2_acc_1877_nl;
  assign Accum2_acc_122_psp_sva_1 = nl_Accum2_acc_122_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1 = (Accum2_acc_123_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[939:935]));
  assign Product1_3_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1259:1255]));
  assign Product1_4_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1579:1575]));
  assign Product1_5_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1899:1895]));
  assign Product1_6_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1890_nl = conv_s2s_11_12(Product1_3_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1890_nl = nl_Accum2_acc_1890_nl[11:0];
  assign nl_Product1_15_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4779:4775]));
  assign Product1_15_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1879_nl = Product1_15_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[299:295]);
  assign Accum2_acc_1879_nl = nl_Accum2_acc_1879_nl[10:0];
  assign nl_Product1_16_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5099:5095]));
  assign Product1_16_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[299:295]));
  assign Product1_1_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[619:615]));
  assign Product1_2_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1893_nl = Accum2_acc_1890_nl + conv_s2s_11_12(Accum2_acc_1879_nl)
      + conv_s2s_11_12(Product1_16_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1893_nl = nl_Accum2_acc_1893_nl[11:0];
  assign nl_Product1_11_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3499:3495]));
  assign Product1_11_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3819:3815]));
  assign Product1_12_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4139:4135]));
  assign Product1_13_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4459:4455]));
  assign Product1_14_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1888_nl = conv_s2s_11_12(Product1_11_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1888_nl = nl_Accum2_acc_1888_nl[11:0];
  assign nl_Product1_7_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2219:2215]));
  assign Product1_7_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2539:2535]));
  assign Product1_8_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2859:2855]));
  assign Product1_9_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3179:3175]));
  assign Product1_10_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1892_nl = Accum2_acc_1888_nl + conv_s2s_11_12(Product1_7_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_60_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1892_nl = nl_Accum2_acc_1892_nl[11:0];
  assign nl_Accum2_acc_123_psp_sva_1 = Accum2_acc_1893_nl + Accum2_acc_1892_nl;
  assign Accum2_acc_123_psp_sva_1 = nl_Accum2_acc_123_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1 = (Accum2_acc_124_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[944:940]));
  assign Product1_3_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1264:1260]));
  assign Product1_4_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1584:1580]));
  assign Product1_5_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1904:1900]));
  assign Product1_6_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1905_nl = conv_s2s_11_12(Product1_3_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1905_nl = nl_Accum2_acc_1905_nl[11:0];
  assign nl_Product1_15_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4784:4780]));
  assign Product1_15_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1894_nl = Product1_15_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[304:300]);
  assign Accum2_acc_1894_nl = nl_Accum2_acc_1894_nl[10:0];
  assign nl_Product1_16_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5104:5100]));
  assign Product1_16_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[304:300]));
  assign Product1_1_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[624:620]));
  assign Product1_2_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1908_nl = Accum2_acc_1905_nl + conv_s2s_11_12(Accum2_acc_1894_nl)
      + conv_s2s_11_12(Product1_16_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1908_nl = nl_Accum2_acc_1908_nl[11:0];
  assign nl_Product1_11_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3504:3500]));
  assign Product1_11_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3824:3820]));
  assign Product1_12_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4144:4140]));
  assign Product1_13_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4464:4460]));
  assign Product1_14_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1903_nl = conv_s2s_11_12(Product1_11_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1903_nl = nl_Accum2_acc_1903_nl[11:0];
  assign nl_Product1_7_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2224:2220]));
  assign Product1_7_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2544:2540]));
  assign Product1_8_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2864:2860]));
  assign Product1_9_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3184:3180]));
  assign Product1_10_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1907_nl = Accum2_acc_1903_nl + conv_s2s_11_12(Product1_7_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_61_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1907_nl = nl_Accum2_acc_1907_nl[11:0];
  assign nl_Accum2_acc_124_psp_sva_1 = Accum2_acc_1908_nl + Accum2_acc_1907_nl;
  assign Accum2_acc_124_psp_sva_1 = nl_Accum2_acc_124_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1 = (Accum2_acc_125_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[949:945]));
  assign Product1_3_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1269:1265]));
  assign Product1_4_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1589:1585]));
  assign Product1_5_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1909:1905]));
  assign Product1_6_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1920_nl = conv_s2s_11_12(Product1_3_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1920_nl = nl_Accum2_acc_1920_nl[11:0];
  assign nl_Product1_15_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4789:4785]));
  assign Product1_15_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1909_nl = Product1_15_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[309:305]);
  assign Accum2_acc_1909_nl = nl_Accum2_acc_1909_nl[10:0];
  assign nl_Product1_16_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5109:5105]));
  assign Product1_16_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[309:305]));
  assign Product1_1_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[629:625]));
  assign Product1_2_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1923_nl = Accum2_acc_1920_nl + conv_s2s_11_12(Accum2_acc_1909_nl)
      + conv_s2s_11_12(Product1_16_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1923_nl = nl_Accum2_acc_1923_nl[11:0];
  assign nl_Product1_11_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3509:3505]));
  assign Product1_11_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3829:3825]));
  assign Product1_12_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4149:4145]));
  assign Product1_13_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4469:4465]));
  assign Product1_14_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1918_nl = conv_s2s_11_12(Product1_11_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1918_nl = nl_Accum2_acc_1918_nl[11:0];
  assign nl_Product1_7_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2229:2225]));
  assign Product1_7_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2549:2545]));
  assign Product1_8_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2869:2865]));
  assign Product1_9_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3189:3185]));
  assign Product1_10_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1922_nl = Accum2_acc_1918_nl + conv_s2s_11_12(Product1_7_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_62_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1922_nl = nl_Accum2_acc_1922_nl[11:0];
  assign nl_Accum2_acc_125_psp_sva_1 = Accum2_acc_1923_nl + Accum2_acc_1922_nl;
  assign Accum2_acc_125_psp_sva_1 = nl_Accum2_acc_125_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1 = (Accum2_acc_126_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[954:950]));
  assign Product1_3_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1274:1270]));
  assign Product1_4_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1594:1590]));
  assign Product1_5_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1914:1910]));
  assign Product1_6_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1935_nl = conv_s2s_11_12(Product1_3_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1935_nl = nl_Accum2_acc_1935_nl[11:0];
  assign nl_Product1_15_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4794:4790]));
  assign Product1_15_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1924_nl = Product1_15_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[314:310]);
  assign Accum2_acc_1924_nl = nl_Accum2_acc_1924_nl[10:0];
  assign nl_Product1_16_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5114:5110]));
  assign Product1_16_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[314:310]));
  assign Product1_1_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[634:630]));
  assign Product1_2_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1938_nl = Accum2_acc_1935_nl + conv_s2s_11_12(Accum2_acc_1924_nl)
      + conv_s2s_11_12(Product1_16_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1938_nl = nl_Accum2_acc_1938_nl[11:0];
  assign nl_Product1_11_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3514:3510]));
  assign Product1_11_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3834:3830]));
  assign Product1_12_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4154:4150]));
  assign Product1_13_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4474:4470]));
  assign Product1_14_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1933_nl = conv_s2s_11_12(Product1_11_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1933_nl = nl_Accum2_acc_1933_nl[11:0];
  assign nl_Product1_7_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2234:2230]));
  assign Product1_7_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2554:2550]));
  assign Product1_8_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2874:2870]));
  assign Product1_9_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3194:3190]));
  assign Product1_10_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1937_nl = Accum2_acc_1933_nl + conv_s2s_11_12(Product1_7_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_63_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1937_nl = nl_Accum2_acc_1937_nl[11:0];
  assign nl_Accum2_acc_126_psp_sva_1 = Accum2_acc_1938_nl + Accum2_acc_1937_nl;
  assign Accum2_acc_126_psp_sva_1 = nl_Accum2_acc_126_psp_sva_1[11:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 = (Accum2_acc_127_psp_sva_1[10:4]!=7'b0000000);
  assign nl_Product1_3_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[17:12])) * $signed((w2_rsci_idat[959:955]));
  assign Product1_3_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_3_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_4_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[23:18])) * $signed((w2_rsci_idat[1279:1275]));
  assign Product1_4_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_4_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_5_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[29:24])) * $signed((w2_rsci_idat[1599:1595]));
  assign Product1_5_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_5_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_6_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[35:30])) * $signed((w2_rsci_idat[1919:1915]));
  assign Product1_6_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_6_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1950_nl = conv_s2s_11_12(Product1_3_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_4_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_5_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_6_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1950_nl = nl_Accum2_acc_1950_nl[11:0];
  assign nl_Product1_15_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[89:84])) * $signed((w2_rsci_idat[4799:4795]));
  assign Product1_15_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_15_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1939_nl = Product1_15_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      + conv_s2s_5_11(b2_rsci_idat[319:315]);
  assign Accum2_acc_1939_nl = nl_Accum2_acc_1939_nl[10:0];
  assign nl_Product1_16_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[95:90])) * $signed((w2_rsci_idat[5119:5115]));
  assign Product1_16_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_16_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_1_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[5:0])) * $signed((w2_rsci_idat[319:315]));
  assign Product1_1_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_1_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_2_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[11:6])) * $signed((w2_rsci_idat[639:635]));
  assign Product1_2_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_2_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1953_nl = Accum2_acc_1950_nl + conv_s2s_11_12(Accum2_acc_1939_nl)
      + conv_s2s_11_12(Product1_16_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_1_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_2_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1953_nl = nl_Accum2_acc_1953_nl[11:0];
  assign nl_Product1_11_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[65:60])) * $signed((w2_rsci_idat[3519:3515]));
  assign Product1_11_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_11_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_12_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[71:66])) * $signed((w2_rsci_idat[3839:3835]));
  assign Product1_12_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_12_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_13_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[77:72])) * $signed((w2_rsci_idat[4159:4155]));
  assign Product1_13_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_13_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_14_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[83:78])) * $signed((w2_rsci_idat[4479:4475]));
  assign Product1_14_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_14_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1948_nl = conv_s2s_11_12(Product1_11_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_12_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_13_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_14_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1948_nl = nl_Accum2_acc_1948_nl[11:0];
  assign nl_Product1_7_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[41:36])) * $signed((w2_rsci_idat[2239:2235]));
  assign Product1_7_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_7_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_8_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[47:42])) * $signed((w2_rsci_idat[2559:2555]));
  assign Product1_8_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_8_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_9_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[53:48])) * $signed((w2_rsci_idat[2879:2875]));
  assign Product1_9_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl =
      nl_Product1_9_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Product1_10_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = $signed(conv_u2s_6_7(input_1_rsci_idat[59:54])) * $signed((w2_rsci_idat[3199:3195]));
  assign Product1_10_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl
      = nl_Product1_10_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl[10:0];
  assign nl_Accum2_acc_1952_nl = Accum2_acc_1948_nl + conv_s2s_11_12(Product1_7_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_8_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_9_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl)
      + conv_s2s_11_12(Product1_10_Product2_64_operator_5_1_true_AC_TRN_AC_WRAP_6_false_mul_nl);
  assign Accum2_acc_1952_nl = nl_Accum2_acc_1952_nl[11:0];
  assign nl_Accum2_acc_127_psp_sva_1 = Accum2_acc_1953_nl + Accum2_acc_1952_nl;
  assign Accum2_acc_127_psp_sva_1 = nl_Accum2_acc_127_psp_sva_1[11:0];
  assign nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[744:740]));
  assign Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[699:695]));
  assign Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[714:710]));
  assign Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[669:665]));
  assign Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[384:380]));
  assign Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[399:395]));
  assign Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[414:410]));
  assign Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[429:425]));
  assign Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[444:440]));
  assign Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[459:455]));
  assign Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[474:470]));
  assign Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[489:485]));
  assign Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[204:200]));
  assign Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[219:215]));
  assign Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[144:140]));
  assign Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[159:155]));
  assign Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[174:170]));
  assign Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[189:185]));
  assign Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[234:230]));
  assign Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[249:245]));
  assign Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[324:320]));
  assign Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[339:335]));
  assign Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[264:260]));
  assign Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[279:275]));
  assign Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[294:290]));
  assign Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[309:305]));
  assign Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[354:350]));
  assign Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[369:365]));
  assign Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[939:935]));
  assign Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[954:950]));
  assign Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[909:905]));
  assign Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[624:620]));
  assign Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[639:635]));
  assign Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[924:920]));
  assign Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[879:875]));
  assign Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[894:890]));
  assign Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[849:845]));
  assign Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[804:800]));
  assign Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[759:755]));
  assign Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[774:770]));
  assign Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[729:725]));
  assign Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[864:860]));
  assign Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[819:815]));
  assign Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[834:830]));
  assign Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[789:785]));
  assign Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_192_nl = conv_s2s_5_6(b5_rsci_idat[9:5]) + conv_s2s_5_6(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[8:4]);
  assign Accum2_1_acc_192_nl = nl_Accum2_1_acc_192_nl[5:0];
  assign nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[684:680]));
  assign Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[654:650]));
  assign Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[84:80]));
  assign Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[99:95]));
  assign Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[114:110]));
  assign Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[129:125]));
  assign Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[24:20]));
  assign Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[39:35]));
  assign Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[54:50]));
  assign Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[69:65]));
  assign Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[564:560]));
  assign Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[579:575]));
  assign Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[594:590]));
  assign Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[609:605]));
  assign Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[504:500]));
  assign Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[519:515]));
  assign Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[534:530]));
  assign Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[549:545]));
  assign Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1 = conv_s2s_9_16(readslicef_15_9_6(Product1_1_50_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_47_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_48_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_45_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_26_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_27_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_28_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_29_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_30_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_31_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_32_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_33_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_14_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_15_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_10_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_11_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_12_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_13_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_16_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_17_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_22_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_23_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_18_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_19_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_20_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_21_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_24_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_25_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_63_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_64_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_61_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_42_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_43_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_62_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_59_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_60_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_57_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_54_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_51_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_52_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_49_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_58_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_55_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_56_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_53_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_10_16({Accum2_1_acc_192_nl , (Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[3:0])})
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_46_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_44_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_6_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_7_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_8_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_9_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_2_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_3_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_4_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_5_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_38_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_39_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_40_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_41_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_34_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_35_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_36_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_37_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1 = nl_Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1[15:0];
  assign nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[719:715]));
  assign Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[734:730]));
  assign Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[689:685]));
  assign Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[704:700]));
  assign Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[374:370]));
  assign Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[389:385]));
  assign Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[404:400]));
  assign Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[419:415]));
  assign Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[434:430]));
  assign Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[449:445]));
  assign Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[464:460]));
  assign Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[479:475]));
  assign Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[194:190]));
  assign Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[209:205]));
  assign Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[134:130]));
  assign Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[149:145]));
  assign Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[164:160]));
  assign Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[179:175]));
  assign Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[224:220]));
  assign Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[239:235]));
  assign Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[314:310]));
  assign Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[329:325]));
  assign Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[254:250]));
  assign Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[269:265]));
  assign Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[284:280]));
  assign Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[299:295]));
  assign Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[344:340]));
  assign Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[359:355]));
  assign Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[929:925]));
  assign Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[944:940]));
  assign Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[959:955]));
  assign Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[614:610]));
  assign Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[629:625]));
  assign Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[899:895]));
  assign Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[914:910]));
  assign Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[869:865]));
  assign Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[884:880]));
  assign Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[779:775]));
  assign Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[794:790]));
  assign Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[749:745]));
  assign Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[764:760]));
  assign Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[839:835]));
  assign Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[854:850]));
  assign Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[809:805]));
  assign Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[824:820]));
  assign Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_193_nl = conv_s2s_5_6(Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[8:4])
      + conv_s2s_5_6(b5_rsci_idat[14:10]);
  assign Accum2_1_acc_193_nl = nl_Accum2_1_acc_193_nl[5:0];
  assign nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[659:655]));
  assign Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[674:670]));
  assign Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[74:70]));
  assign Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[89:85]));
  assign Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[104:100]));
  assign Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[119:115]));
  assign Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_4_9 , layer4_out_conc_4_8_6 , ({{3{layer4_out_0_2_lpi_1_dfm_1}},
      layer4_out_0_2_lpi_1_dfm_1}) , layer4_out_0_2_lpi_1_dfm_1 , layer4_out_0_2_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[14:10]));
  assign Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[29:25]));
  assign Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[44:40]));
  assign Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[59:55]));
  assign Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[554:550]));
  assign Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[569:565]));
  assign Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[584:580]));
  assign Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[599:595]));
  assign Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[494:490]));
  assign Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[509:505]));
  assign Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[524:520]));
  assign Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[539:535]));
  assign Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1 = conv_s2s_9_16(readslicef_15_9_6(Product1_1_48_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_49_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_46_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_47_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_25_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_26_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_27_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_28_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_29_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_30_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_31_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_32_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_13_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_14_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_9_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_10_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_11_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_12_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_15_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_16_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_21_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_22_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_17_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_18_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_19_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_20_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_23_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_24_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_62_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_63_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_64_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_41_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_42_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_60_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_61_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_58_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_59_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_52_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_53_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_50_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_51_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_56_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_57_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_54_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_55_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_10_16({Accum2_1_acc_193_nl , (Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[3:0])})
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_44_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_45_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_5_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_6_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_7_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_8_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_1_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_2_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_3_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_4_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_37_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_38_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_39_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_40_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_33_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_34_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_35_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_36_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1 = nl_Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1[15:0];
  assign nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[739:735]));
  assign Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[694:690]));
  assign Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[709:705]));
  assign Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[664:660]));
  assign Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[379:375]));
  assign Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[394:390]));
  assign Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[409:405]));
  assign Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[424:420]));
  assign Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[439:435]));
  assign Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[454:450]));
  assign Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[469:465]));
  assign Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[484:480]));
  assign Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[199:195]));
  assign Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[214:210]));
  assign Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[139:135]));
  assign Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[154:150]));
  assign Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[169:165]));
  assign Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[184:180]));
  assign Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[229:225]));
  assign Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[244:240]));
  assign Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[319:315]));
  assign Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[334:330]));
  assign Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[259:255]));
  assign Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[274:270]));
  assign Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[289:285]));
  assign Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[304:300]));
  assign Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[349:345]));
  assign Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[364:360]));
  assign Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[934:930]));
  assign Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[949:945]));
  assign Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[904:900]));
  assign Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[619:615]));
  assign Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[634:630]));
  assign Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[919:915]));
  assign Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[874:870]));
  assign Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[889:885]));
  assign Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[844:840]));
  assign Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[799:795]));
  assign Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[754:750]));
  assign Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[769:765]));
  assign Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[724:720]));
  assign Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[859:855]));
  assign Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[814:810]));
  assign Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[829:825]));
  assign Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[784:780]));
  assign Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum2_1_acc_191_nl = conv_s2s_5_6(b5_rsci_idat[4:0]) + conv_s2s_5_6(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[8:4]);
  assign Accum2_1_acc_191_nl = nl_Accum2_1_acc_191_nl[5:0];
  assign nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[679:675]));
  assign Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[649:645]));
  assign Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[79:75]));
  assign Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[94:90]));
  assign Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[109:105]));
  assign Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[124:120]));
  assign Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[19:15]));
  assign Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[34:30]));
  assign Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[49:45]));
  assign Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[64:60]));
  assign Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[559:555]));
  assign Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[574:570]));
  assign Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[589:585]));
  assign Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[604:600]));
  assign Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[499:495]));
  assign Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[514:510]));
  assign Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[529:525]));
  assign Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[544:540]));
  assign Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign nl_Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1 = conv_s2s_9_16(readslicef_15_9_6(Product1_1_50_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_47_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_48_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_45_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_26_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_27_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_28_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_29_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_30_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_31_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_32_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_33_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_14_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_15_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_10_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_11_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_12_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_13_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_16_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_17_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_22_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_23_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_18_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_19_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_20_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_21_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_24_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_25_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_63_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_64_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_61_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_42_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_43_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_62_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_59_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_60_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_57_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_54_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_51_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_52_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_49_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_58_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_55_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_56_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_53_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_10_16({Accum2_1_acc_191_nl , (Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1[3:0])})
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_46_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_44_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_6_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_7_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_8_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_9_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_2_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_3_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_4_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_5_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_38_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_39_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_40_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_41_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_34_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_35_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_36_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl))
      + conv_s2s_9_16(readslicef_15_9_6(Product1_1_37_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl));
  assign Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1 = nl_Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1[15:0];
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_12_1;
  assign nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_6 , ({{3{nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1}},
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1})
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1
      , nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[644:640]));
  assign Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1
      = readslicef_15_9_6(Product1_1_43_Product2_1_3_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign layer4_out_0_2_lpi_1_dfm_1 = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1
      & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_conc_13_pmx_1_lpi_1_dfm_1
      = nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1 & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_12_1;
  assign nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_4_9 , layer4_out_conc_4_8_6 , ({{3{layer4_out_0_2_lpi_1_dfm_1}},
      layer4_out_0_2_lpi_1_dfm_1}) , layer4_out_0_2_lpi_1_dfm_1 , layer4_out_0_2_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[9:5]));
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1
      = readslicef_15_9_6(Product1_1_1_Product2_1_2_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = $signed(conv_u2s_10_11({layer4_out_conc_4_9 , layer4_out_conc_4_8_6 , ({{3{layer4_out_0_2_lpi_1_dfm_1}},
      layer4_out_0_2_lpi_1_dfm_1}) , layer4_out_0_2_lpi_1_dfm_1 , layer4_out_0_2_lpi_1_dfm_1}))
      * $signed((w5_rsci_idat[4:0]));
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl
      = nl_Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl[14:0];
  assign Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_itm_14_6_1
      = readslicef_15_9_6(Product1_1_1_Product2_1_1_nnet_product_mult_layer4_t_config6_weight_t_product_mul_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl =  -conv_s2s_12_13(Accum2_acc_127_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl =  -conv_s2s_12_13(Accum2_acc_126_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl =  -conv_s2s_12_13(Accum2_acc_125_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl =  -conv_s2s_12_13(Accum2_acc_124_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl =  -conv_s2s_12_13(Accum2_acc_123_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl =  -conv_s2s_12_13(Accum2_acc_122_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl =  -conv_s2s_12_13(Accum2_acc_121_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl =  -conv_s2s_12_13(Accum2_acc_120_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl =  -conv_s2s_12_13(Accum2_acc_119_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl =  -conv_s2s_12_13(Accum2_acc_118_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl =  -conv_s2s_12_13(Accum2_acc_117_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl =  -conv_s2s_12_13(Accum2_acc_116_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl =  -conv_s2s_12_13(Accum2_acc_115_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl =  -conv_s2s_12_13(Accum2_acc_114_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl =  -conv_s2s_12_13(Accum2_acc_113_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl =  -conv_s2s_12_13(Accum2_acc_112_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl =  -conv_s2s_12_13(Accum2_acc_111_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl =  -conv_s2s_12_13(Accum2_acc_110_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl =  -conv_s2s_12_13(Accum2_acc_109_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl =  -conv_s2s_12_13(Accum2_acc_108_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl =  -conv_s2s_12_13(Accum2_acc_107_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl =  -conv_s2s_12_13(Accum2_acc_106_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl =  -conv_s2s_12_13(Accum2_acc_105_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl =  -conv_s2s_12_13(Accum2_acc_104_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl =  -conv_s2s_12_13(Accum2_acc_103_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl =  -conv_s2s_12_13(Accum2_acc_102_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl =  -conv_s2s_12_13(Accum2_acc_101_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl =  -conv_s2s_12_13(Accum2_acc_100_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl =  -conv_s2s_12_13(Accum2_acc_99_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl =  -conv_s2s_12_13(Accum2_acc_98_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl =  -conv_s2s_12_13(Accum2_acc_97_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl =  -conv_s2s_12_13(Accum2_acc_96_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl =  -conv_s2s_12_13(Accum2_acc_95_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl =  -conv_s2s_12_13(Accum2_acc_94_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl =  -conv_s2s_12_13(Accum2_acc_93_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl =  -conv_s2s_12_13(Accum2_acc_92_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl =  -conv_s2s_12_13(Accum2_acc_91_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl =  -conv_s2s_12_13(Accum2_acc_90_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl =  -conv_s2s_12_13(Accum2_acc_89_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl =  -conv_s2s_12_13(Accum2_acc_88_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl =  -conv_s2s_12_13(Accum2_acc_87_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl =  -conv_s2s_12_13(Accum2_acc_86_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl =  -conv_s2s_12_13(Accum2_acc_85_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl =  -conv_s2s_12_13(Accum2_acc_84_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl =  -conv_s2s_12_13(Accum2_acc_83_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl =  -conv_s2s_12_13(Accum2_acc_82_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl =  -conv_s2s_12_13(Accum2_acc_81_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl =  -conv_s2s_12_13(Accum2_acc_80_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl =  -conv_s2s_12_13(Accum2_acc_79_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl =  -conv_s2s_12_13(Accum2_acc_78_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl =  -conv_s2s_12_13(Accum2_acc_77_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl =  -conv_s2s_12_13(Accum2_acc_76_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl =  -conv_s2s_12_13(Accum2_acc_75_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl =  -conv_s2s_12_13(Accum2_acc_74_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl =  -conv_s2s_12_13(Accum2_acc_73_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl =  -conv_s2s_12_13(Accum2_acc_72_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl =  -conv_s2s_12_13(Accum2_acc_71_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl =  -conv_s2s_12_13(Accum2_acc_70_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl =  -conv_s2s_12_13(Accum2_acc_69_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl =  -conv_s2s_12_13(Accum2_acc_68_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl =  -conv_s2s_12_13(Accum2_acc_67_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl =  -conv_s2s_12_13(Accum2_acc_66_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl =  -conv_s2s_12_13(Accum2_acc_65_psp_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_nl);
  assign nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl =  -conv_s2s_12_13(layer3_out_0_15_4_sva_1);
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl = nl_operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl[12:0];
  assign operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_12_1 = readslicef_13_1_12(operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_nl);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_9 = ((Accum2_acc_104_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_104_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_41_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_204_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_41_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_39_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_9 = ((Accum2_acc_105_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_105_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_42_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_206_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_42_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_40_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_9 = ((Accum2_acc_125_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_125_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_62_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_208_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_62_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_60_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_9 = ((Accum2_acc_126_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_126_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_63_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_210_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_63_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_61_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_9 = ((Accum2_acc_127_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_127_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_212_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_64_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_62_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_9 = ((Accum2_acc_123_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_123_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_60_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_214_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_60_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_58_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_9 = ((Accum2_acc_124_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_124_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_61_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_216_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_61_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_59_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_9 = ((Accum2_acc_121_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_121_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_58_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_218_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_58_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_56_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_9 = ((Accum2_acc_122_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_122_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_59_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_220_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_59_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_57_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_9 = ((Accum2_acc_119_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_119_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_56_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_222_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_56_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_54_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_9 = ((Accum2_acc_120_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_120_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_57_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_224_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_57_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_55_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_9 = ((Accum2_acc_117_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_117_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_54_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_226_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_54_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_52_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_9 = ((Accum2_acc_118_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_118_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_55_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_228_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_55_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_53_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_9 = ((Accum2_acc_115_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_115_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_52_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_230_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_52_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_50_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_9 = ((Accum2_acc_116_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_116_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_53_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_232_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_53_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_51_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_9 = ((Accum2_acc_113_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_113_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_50_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_234_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_50_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_48_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_9 = ((Accum2_acc_114_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_114_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_51_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_236_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_51_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_49_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_9 = ((Accum2_acc_111_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_111_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_48_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_238_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_48_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_46_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_9 = ((Accum2_acc_112_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_112_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_49_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_240_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_49_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_47_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_9 = ((Accum2_acc_109_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_109_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_46_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_242_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_46_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_44_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_9 = ((Accum2_acc_110_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_110_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_47_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_244_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_47_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_45_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_9 = ((Accum2_acc_107_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_107_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_44_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_246_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_44_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_42_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_9 = ((Accum2_acc_108_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_108_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_45_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_248_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_45_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_43_itm_12_1);
  assign layer4_out_conc_4_9 = ((layer3_out_0_15_4_sva_1[3]) | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1)
      & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((layer3_out_0_15_4_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_1_sva_1);
  assign layer4_out_conc_4_8_6 = MUX_v_3_2_2(3'b000, nnet_relu_layer3_t_layer4_t_relu_config4_for_1_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_63_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_9 = ((Accum2_acc_65_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_65_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_2_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_250_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_2_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_9 = ((Accum2_acc_66_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_66_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_3_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_252_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_3_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_1_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_9 = ((Accum2_acc_67_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_67_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_4_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_254_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_4_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_2_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_9 = ((Accum2_acc_68_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_68_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_5_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_256_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_5_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_3_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_9 = ((Accum2_acc_69_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_69_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_6_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_258_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_6_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_4_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_9 = ((Accum2_acc_70_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_70_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_7_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_260_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_7_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_5_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_9 = ((Accum2_acc_71_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_71_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_8_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_262_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_8_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_6_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_9 = ((Accum2_acc_72_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_72_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_9_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_264_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_9_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_7_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_9 = ((Accum2_acc_73_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_73_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_10_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_266_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_10_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_8_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_9 = ((Accum2_acc_74_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_74_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_11_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_268_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_11_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_9_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_9 = ((Accum2_acc_75_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_75_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_12_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_270_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_12_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_10_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_9 = ((Accum2_acc_76_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_76_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_13_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_272_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_13_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_11_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_9 = ((Accum2_acc_77_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_77_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_14_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_274_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_14_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_12_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_9 = ((Accum2_acc_78_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_78_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_15_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_276_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_15_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_13_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_9 = ((Accum2_acc_79_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_79_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_16_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_278_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_16_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_14_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_9 = ((Accum2_acc_80_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_80_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_17_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_280_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_17_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_15_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_9 = ((Accum2_acc_81_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_81_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_18_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_282_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_18_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_16_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_9 = ((Accum2_acc_82_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_82_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_19_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_284_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_19_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_17_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_9 = ((Accum2_acc_83_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_83_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_20_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_286_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_20_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_18_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_9 = ((Accum2_acc_84_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_84_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_21_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_288_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_21_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_19_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_9 = ((Accum2_acc_85_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_85_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_22_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_290_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_22_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_20_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_9 = ((Accum2_acc_86_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_86_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_23_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_292_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_23_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_21_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_9 = ((Accum2_acc_87_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_87_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_24_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_294_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_24_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_22_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_9 = ((Accum2_acc_88_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_88_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_25_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_296_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_25_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_23_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_9 = ((Accum2_acc_89_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_89_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_26_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_298_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_26_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_24_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_9 = ((Accum2_acc_90_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_90_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_27_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_300_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_27_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_25_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_9 = ((Accum2_acc_91_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_91_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_28_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_302_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_28_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_26_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_9 = ((Accum2_acc_92_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_92_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_29_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_304_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_29_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_27_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_9 = ((Accum2_acc_93_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_93_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_30_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_306_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_30_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_28_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_9 = ((Accum2_acc_94_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_94_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_31_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_308_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_31_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_29_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_9 = ((Accum2_acc_95_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_95_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_32_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_310_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_32_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_30_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_9 = ((Accum2_acc_96_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_96_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_33_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_312_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_33_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_31_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_9 = ((Accum2_acc_97_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_97_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_34_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_314_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_34_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_32_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_9 = ((Accum2_acc_98_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_98_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_35_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_316_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_35_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_33_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_9 = ((Accum2_acc_99_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_99_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_36_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_318_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_36_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_34_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_9 = ((Accum2_acc_100_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_100_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_37_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_320_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_37_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_35_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_9 = ((Accum2_acc_101_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_101_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_38_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_322_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_38_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_36_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_9 = ((Accum2_acc_102_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_102_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_39_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_324_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_39_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_37_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_9 = ((Accum2_acc_103_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_103_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_40_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_326_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_40_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_38_itm_12_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_9 = ((Accum2_acc_106_psp_sva_1[3])
      | nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1) & operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_12_1;
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl
      = MUX_v_3_2_2((Accum2_acc_106_psp_sva_1[2:0]), 3'b111, nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nor_ovfl_43_sva_1);
  assign nnet_relu_layer3_t_layer4_t_relu_config4_for_if_conc_328_8_6 = MUX_v_3_2_2(3'b000,
      nnet_relu_layer3_t_layer4_t_relu_config4_for_43_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_nnet_relu_layer3_t_layer4_t_relu_config4_for_if_or_2_nl,
      operator_16_8_true_AC_RND_CONV_AC_SAT_acc_41_itm_12_1);
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat <= 2'b00;
    end
    else begin
      layer7_out_rsci_idat <= ~(MUX_v_2_2_2(argmax_else_mux_nl, 2'b11, argmax_if_argmax_if_argmax_if_nor_nl));
    end
  end
  assign nl_argmax_else_aif_acc_nl = Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1
      - Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1;
  assign argmax_else_aif_acc_nl = nl_argmax_else_aif_acc_nl[15:0];
  assign nl_argmax_else_acc_nl = Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1
      - Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1;
  assign argmax_else_acc_nl = nl_argmax_else_acc_nl[15:0];
  assign argmax_else_if_argmax_else_if_argmax_else_if_nor_nl = ~((readslicef_16_1_15(argmax_else_aif_acc_nl))
      | (readslicef_16_1_15(argmax_else_acc_nl)));
  assign argmax_else_mux_nl = MUX_v_2_2_2(2'b01, 2'b10, argmax_else_if_argmax_else_if_argmax_else_if_nor_nl);
  assign nl_argmax_aif_acc_nl = Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1
      - Accum1_1_64_Accum2_1_3_Accum2_1_acc_1_ncse_sva_1;
  assign argmax_aif_acc_nl = nl_argmax_aif_acc_nl[15:0];
  assign nl_argmax_acc_nl = Accum1_1_64_Accum2_1_1_Accum2_1_acc_1_ncse_sva_1 - Accum1_1_64_Accum2_1_2_Accum2_1_acc_1_ncse_sva_1;
  assign argmax_acc_nl = nl_argmax_acc_nl[15:0];
  assign argmax_if_argmax_if_argmax_if_nor_nl = ~((readslicef_16_1_15(argmax_aif_acc_nl))
      | (readslicef_16_1_15(argmax_acc_nl)));

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [8:0] readslicef_15_9_6;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_15_9_6 = tmp[8:0];
  end
  endfunction


  function automatic [0:0] readslicef_16_1_15;
    input [15:0] vector;
    reg [15:0] tmp;
  begin
    tmp = vector >> 15;
    readslicef_16_1_15 = tmp[0:0];
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_5_11 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_11 = {{6{vector[4]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_9_16 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_16 = {{7{vector[8]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_10_16 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_16 = {{6{vector[9]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    myproject
// ------------------------------------------------------------------


module myproject (
  clk, rst, input_1_rsc_dat, layer7_out_rsc_dat, w2_rsc_dat, b2_rsc_dat, w5_rsc_dat,
      b5_rsc_dat
);
  input clk;
  input rst;
  input [95:0] input_1_rsc_dat;
  output [1:0] layer7_out_rsc_dat;
  input [5119:0] w2_rsc_dat;
  input [319:0] b2_rsc_dat;
  input [959:0] w5_rsc_dat;
  input [14:0] b5_rsc_dat;



  // Interconnect Declarations for Component Instantiations 
  converterBlock_myproject_core myproject_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .w2_rsc_dat(w2_rsc_dat),
      .b2_rsc_dat(b2_rsc_dat),
      .w5_rsc_dat(w5_rsc_dat),
      .b5_rsc_dat(b5_rsc_dat)
    );
endmodule



